
module Homework3_3_LUT_interpolation(clk,in_theta,realout,imagout);
input [11:0]in_theta;
input clk;
output [15:0]realout;
output [15:0]imagout;


wire [11:0]in_theta;
wire clk;
reg [15:0]realout;
reg [15:0]imagout;

reg [11:0]theta;
reg [11:0]thegen1;
reg [11:0]thegen;
reg [15:0]real3;
reg [15:0]imag3;
reg [15:0]real2;
reg [15:0]imag2;
reg [15:0]real1;
reg [15:0]imag1;
reg [15:0]tmp;
reg [15:0]tmpreal1;
reg [15:0]tmpreal2;
reg [15:0]tmpimag1;
reg [15:0]tmpimag2;


always@(posedge clk)begin
theta<= #1 in_theta;
realout<=#1 real3;
imagout<=#1 imag3;
end

always @(*) begin
if (theta<=12'b010000000000)begin
	thegen = theta;
	real3=real2;
	imag3=imag2;
	end
else if (theta<=12'b100000000000 && theta>12'b010000000000)begin
	thegen = 12'b100000000000-theta;
	real3 =~real2+1'b1;
	imag3=imag2;
	end
else if (theta<=12'b110000000000 && theta>12'b100000000000)begin
	thegen = theta-12'b100000000000;
	real3 =~real2+1'b1;
	imag3=~imag2+1'b1;
	end
else if (theta<=12'b111111111111 && theta>12'b110000000000)begin
	thegen = 12'b111111111111-theta+1'b1;
	real3 =real2;
	imag3=~imag2+1'b1;
	end

if (thegen>12'b001000000000 && thegen[0]== 1'b0)begin
	thegen1=12'b010000000000-thegen;
	tmp=imag1;	
	imag2=real1;	
	real2=tmp;
end
else if(thegen<=12'b001000000000 && thegen[0]==1'b0)begin
	thegen1=thegen;
	imag2=imag1;	
	real2=real1;
end
else if (thegen>12'b001000000000 && thegen[0]==1'b1)begin
	thegen=12'b010000000010-thegen;
	thegen1=thegen+1'b1;
	tmpreal1=real1;
	tmpimag1=imag1;
	thegen1=#1 thegen-1'b1;
	tmpreal2= real1;
	tmpimag2= imag1;
	imag2=({tmpimag2[15],tmpimag2[15],tmpimag2[15],tmpimag2}+{tmpimag1[15],tmpimag1[15],tmpimag1[15],tmpimag1}+1'b1)>>1;
	real2=({tmpreal2[15],tmpreal2[15],tmpreal2[15],tmpreal2}+{tmpreal1[15],tmpreal1[15],tmpreal1[15],tmpreal1}+1'b1)>>1;
	tmp=imag1;	
	imag2=real1;	
	real2=tmp;
end
else if(thegen<=12'b001000000000 && thegen[0]==1'b1)begin	
	thegen1=thegen+1'b1;
	tmpreal1=real1;
	tmpimag1=imag1;
	thegen1=#3 thegen-1'b1;
	tmpreal2= real1;
	tmpimag2= imag1;
	imag2=({tmpimag2[15],tmpimag2[15],tmpimag2[15],tmpimag2}+{tmpimag1[15],tmpimag1[15],tmpimag1[15],tmpimag1}+1'b1)>>1;
	real2=({tmpreal2[15],tmpreal2[15],tmpreal2[15],tmpreal2}+{tmpreal1[15],tmpreal1[15],tmpreal1[15],tmpreal1}+1'b1)>>1;
	$display(tmpreal1);
	$display(tmpreal2);
	$display(real2);
	$display("-----");
end
end


always @(thegen1) begin
  case (thegen1)
    12'b000000000000: begin  real1=16'b0100000000000000; imag1=16'b0000000000000000;  end  // angle = 0.000000 pi
    12'b000000000010: begin  real1=16'b0100000000000000; imag1=16'b0000000000110010;  end  // angle = 0.000977 pi
    12'b000000000100: begin  real1=16'b0100000000000000; imag1=16'b0000000001100101;  end  // angle = 0.001953 pi
    12'b000000000110: begin  real1=16'b0011111111111111; imag1=16'b0000000010010111;  end  // angle = 0.002930 pi
    12'b000000001000: begin  real1=16'b0011111111111111; imag1=16'b0000000011001001;  end  // angle = 0.003906 pi
    12'b000000001010: begin  real1=16'b0011111111111110; imag1=16'b0000000011111011;  end  // angle = 0.004883 pi
    12'b000000001100: begin  real1=16'b0011111111111101; imag1=16'b0000000100101110;  end  // angle = 0.005859 pi
    12'b000000001110: begin  real1=16'b0011111111111100; imag1=16'b0000000101100000;  end  // angle = 0.006836 pi
    12'b000000010000: begin  real1=16'b0011111111111011; imag1=16'b0000000110010010;  end  // angle = 0.007812 pi
    12'b000000010010: begin  real1=16'b0011111111111010; imag1=16'b0000000111000100;  end  // angle = 0.008789 pi
    12'b000000010100: begin  real1=16'b0011111111111000; imag1=16'b0000000111110111;  end  // angle = 0.009766 pi
    12'b000000010110: begin  real1=16'b0011111111110111; imag1=16'b0000001000101001;  end  // angle = 0.010742 pi
    12'b000000011000: begin  real1=16'b0011111111110101; imag1=16'b0000001001011011;  end  // angle = 0.011719 pi
    12'b000000011010: begin  real1=16'b0011111111110011; imag1=16'b0000001010001101;  end  // angle = 0.012695 pi
    12'b000000011100: begin  real1=16'b0011111111110001; imag1=16'b0000001011000000;  end  // angle = 0.013672 pi
    12'b000000011110: begin  real1=16'b0011111111101111; imag1=16'b0000001011110010;  end  // angle = 0.014648 pi
    12'b000000100000: begin  real1=16'b0011111111101100; imag1=16'b0000001100100100;  end  // angle = 0.015625 pi
    12'b000000100010: begin  real1=16'b0011111111101010; imag1=16'b0000001101010110;  end  // angle = 0.016602 pi
    12'b000000100100: begin  real1=16'b0011111111100111; imag1=16'b0000001110001000;  end  // angle = 0.017578 pi
    12'b000000100110: begin  real1=16'b0011111111100100; imag1=16'b0000001110111011;  end  // angle = 0.018555 pi
    12'b000000101000: begin  real1=16'b0011111111100001; imag1=16'b0000001111101101;  end  // angle = 0.019531 pi
    12'b000000101010: begin  real1=16'b0011111111011110; imag1=16'b0000010000011111;  end  // angle = 0.020508 pi
    12'b000000101100: begin  real1=16'b0011111111011011; imag1=16'b0000010001010001;  end  // angle = 0.021484 pi
    12'b000000101110: begin  real1=16'b0011111111010111; imag1=16'b0000010010000011;  end  // angle = 0.022461 pi
    12'b000000110000: begin  real1=16'b0011111111010100; imag1=16'b0000010010110101;  end  // angle = 0.023438 pi
    12'b000000110010: begin  real1=16'b0011111111010000; imag1=16'b0000010011100111;  end  // angle = 0.024414 pi
    12'b000000110100: begin  real1=16'b0011111111001100; imag1=16'b0000010100011010;  end  // angle = 0.025391 pi
    12'b000000110110: begin  real1=16'b0011111111001000; imag1=16'b0000010101001100;  end  // angle = 0.026367 pi
    12'b000000111000: begin  real1=16'b0011111111000100; imag1=16'b0000010101111110;  end  // angle = 0.027344 pi
    12'b000000111010: begin  real1=16'b0011111110111111; imag1=16'b0000010110110000;  end  // angle = 0.028320 pi
    12'b000000111100: begin  real1=16'b0011111110111011; imag1=16'b0000010111100010;  end  // angle = 0.029297 pi
    12'b000000111110: begin  real1=16'b0011111110110110; imag1=16'b0000011000010100;  end  // angle = 0.030273 pi
    12'b000001000000: begin  real1=16'b0011111110110001; imag1=16'b0000011001000110;  end  // angle = 0.031250 pi
    12'b000001000010: begin  real1=16'b0011111110101100; imag1=16'b0000011001111000;  end  // angle = 0.032227 pi
    12'b000001000100: begin  real1=16'b0011111110100111; imag1=16'b0000011010101010;  end  // angle = 0.033203 pi
    12'b000001000110: begin  real1=16'b0011111110100010; imag1=16'b0000011011011100;  end  // angle = 0.034180 pi
    12'b000001001000: begin  real1=16'b0011111110011100; imag1=16'b0000011100001110;  end  // angle = 0.035156 pi
    12'b000001001010: begin  real1=16'b0011111110010111; imag1=16'b0000011101000000;  end  // angle = 0.036133 pi
    12'b000001001100: begin  real1=16'b0011111110010001; imag1=16'b0000011101110010;  end  // angle = 0.037109 pi
    12'b000001001110: begin  real1=16'b0011111110001011; imag1=16'b0000011110100100;  end  // angle = 0.038086 pi
    12'b000001010000: begin  real1=16'b0011111110000101; imag1=16'b0000011111010110;  end  // angle = 0.039062 pi
    12'b000001010010: begin  real1=16'b0011111101111111; imag1=16'b0000100000000111;  end  // angle = 0.040039 pi
    12'b000001010100: begin  real1=16'b0011111101111000; imag1=16'b0000100000111001;  end  // angle = 0.041016 pi
    12'b000001010110: begin  real1=16'b0011111101110010; imag1=16'b0000100001101011;  end  // angle = 0.041992 pi
    12'b000001011000: begin  real1=16'b0011111101101011; imag1=16'b0000100010011101;  end  // angle = 0.042969 pi
    12'b000001011010: begin  real1=16'b0011111101100100; imag1=16'b0000100011001111;  end  // angle = 0.043945 pi
    12'b000001011100: begin  real1=16'b0011111101011101; imag1=16'b0000100100000001;  end  // angle = 0.044922 pi
    12'b000001011110: begin  real1=16'b0011111101010110; imag1=16'b0000100100110010;  end  // angle = 0.045898 pi
    12'b000001100000: begin  real1=16'b0011111101001111; imag1=16'b0000100101100100;  end  // angle = 0.046875 pi
    12'b000001100010: begin  real1=16'b0011111101000111; imag1=16'b0000100110010110;  end  // angle = 0.047852 pi
    12'b000001100100: begin  real1=16'b0011111101000000; imag1=16'b0000100111000111;  end  // angle = 0.048828 pi
    12'b000001100110: begin  real1=16'b0011111100111000; imag1=16'b0000100111111001;  end  // angle = 0.049805 pi
    12'b000001101000: begin  real1=16'b0011111100110000; imag1=16'b0000101000101011;  end  // angle = 0.050781 pi
    12'b000001101010: begin  real1=16'b0011111100101000; imag1=16'b0000101001011100;  end  // angle = 0.051758 pi
    12'b000001101100: begin  real1=16'b0011111100100000; imag1=16'b0000101010001110;  end  // angle = 0.052734 pi
    12'b000001101110: begin  real1=16'b0011111100010111; imag1=16'b0000101011000000;  end  // angle = 0.053711 pi
    12'b000001110000: begin  real1=16'b0011111100001111; imag1=16'b0000101011110001;  end  // angle = 0.054688 pi
    12'b000001110010: begin  real1=16'b0011111100000110; imag1=16'b0000101100100011;  end  // angle = 0.055664 pi
    12'b000001110100: begin  real1=16'b0011111011111101; imag1=16'b0000101101010100;  end  // angle = 0.056641 pi
    12'b000001110110: begin  real1=16'b0011111011110100; imag1=16'b0000101110000101;  end  // angle = 0.057617 pi
    12'b000001111000: begin  real1=16'b0011111011101011; imag1=16'b0000101110110111;  end  // angle = 0.058594 pi
    12'b000001111010: begin  real1=16'b0011111011100010; imag1=16'b0000101111101000;  end  // angle = 0.059570 pi
    12'b000001111100: begin  real1=16'b0011111011011000; imag1=16'b0000110000011010;  end  // angle = 0.060547 pi
    12'b000001111110: begin  real1=16'b0011111011001111; imag1=16'b0000110001001011;  end  // angle = 0.061523 pi
    12'b000010000000: begin  real1=16'b0011111011000101; imag1=16'b0000110001111100;  end  // angle = 0.062500 pi
    12'b000010000010: begin  real1=16'b0011111010111011; imag1=16'b0000110010101110;  end  // angle = 0.063477 pi
    12'b000010000100: begin  real1=16'b0011111010110001; imag1=16'b0000110011011111;  end  // angle = 0.064453 pi
    12'b000010000110: begin  real1=16'b0011111010100111; imag1=16'b0000110100010000;  end  // angle = 0.065430 pi
    12'b000010001000: begin  real1=16'b0011111010011101; imag1=16'b0000110101000001;  end  // angle = 0.066406 pi
    12'b000010001010: begin  real1=16'b0011111010010010; imag1=16'b0000110101110010;  end  // angle = 0.067383 pi
    12'b000010001100: begin  real1=16'b0011111010001000; imag1=16'b0000110110100100;  end  // angle = 0.068359 pi
    12'b000010001110: begin  real1=16'b0011111001111101; imag1=16'b0000110111010101;  end  // angle = 0.069336 pi
    12'b000010010000: begin  real1=16'b0011111001110010; imag1=16'b0000111000000110;  end  // angle = 0.070312 pi
    12'b000010010010: begin  real1=16'b0011111001100111; imag1=16'b0000111000110111;  end  // angle = 0.071289 pi
    12'b000010010100: begin  real1=16'b0011111001011100; imag1=16'b0000111001101000;  end  // angle = 0.072266 pi
    12'b000010010110: begin  real1=16'b0011111001010000; imag1=16'b0000111010011001;  end  // angle = 0.073242 pi
    12'b000010011000: begin  real1=16'b0011111001000101; imag1=16'b0000111011001010;  end  // angle = 0.074219 pi
    12'b000010011010: begin  real1=16'b0011111000111001; imag1=16'b0000111011111011;  end  // angle = 0.075195 pi
    12'b000010011100: begin  real1=16'b0011111000101101; imag1=16'b0000111100101011;  end  // angle = 0.076172 pi
    12'b000010011110: begin  real1=16'b0011111000100001; imag1=16'b0000111101011100;  end  // angle = 0.077148 pi
    12'b000010100000: begin  real1=16'b0011111000010101; imag1=16'b0000111110001101;  end  // angle = 0.078125 pi
    12'b000010100010: begin  real1=16'b0011111000001001; imag1=16'b0000111110111110;  end  // angle = 0.079102 pi
    12'b000010100100: begin  real1=16'b0011110111111100; imag1=16'b0000111111101110;  end  // angle = 0.080078 pi
    12'b000010100110: begin  real1=16'b0011110111110000; imag1=16'b0001000000011111;  end  // angle = 0.081055 pi
    12'b000010101000: begin  real1=16'b0011110111100011; imag1=16'b0001000001010000;  end  // angle = 0.082031 pi
    12'b000010101010: begin  real1=16'b0011110111010110; imag1=16'b0001000010000000;  end  // angle = 0.083008 pi
    12'b000010101100: begin  real1=16'b0011110111001001; imag1=16'b0001000010110001;  end  // angle = 0.083984 pi
    12'b000010101110: begin  real1=16'b0011110110111100; imag1=16'b0001000011100001;  end  // angle = 0.084961 pi
    12'b000010110000: begin  real1=16'b0011110110101111; imag1=16'b0001000100010010;  end  // angle = 0.085937 pi
    12'b000010110010: begin  real1=16'b0011110110100001; imag1=16'b0001000101000010;  end  // angle = 0.086914 pi
    12'b000010110100: begin  real1=16'b0011110110010011; imag1=16'b0001000101110011;  end  // angle = 0.087891 pi
    12'b000010110110: begin  real1=16'b0011110110000110; imag1=16'b0001000110100011;  end  // angle = 0.088867 pi
    12'b000010111000: begin  real1=16'b0011110101111000; imag1=16'b0001000111010011;  end  // angle = 0.089844 pi
    12'b000010111010: begin  real1=16'b0011110101101010; imag1=16'b0001001000000100;  end  // angle = 0.090820 pi
    12'b000010111100: begin  real1=16'b0011110101011011; imag1=16'b0001001000110100;  end  // angle = 0.091797 pi
    12'b000010111110: begin  real1=16'b0011110101001101; imag1=16'b0001001001100100;  end  // angle = 0.092773 pi
    12'b000011000000: begin  real1=16'b0011110100111111; imag1=16'b0001001010010100;  end  // angle = 0.093750 pi
    12'b000011000010: begin  real1=16'b0011110100110000; imag1=16'b0001001011000100;  end  // angle = 0.094727 pi
    12'b000011000100: begin  real1=16'b0011110100100001; imag1=16'b0001001011110100;  end  // angle = 0.095703 pi
    12'b000011000110: begin  real1=16'b0011110100010010; imag1=16'b0001001100100100;  end  // angle = 0.096680 pi
    12'b000011001000: begin  real1=16'b0011110100000011; imag1=16'b0001001101010100;  end  // angle = 0.097656 pi
    12'b000011001010: begin  real1=16'b0011110011110100; imag1=16'b0001001110000100;  end  // angle = 0.098633 pi
    12'b000011001100: begin  real1=16'b0011110011100100; imag1=16'b0001001110110100;  end  // angle = 0.099609 pi
    12'b000011001110: begin  real1=16'b0011110011010101; imag1=16'b0001001111100100;  end  // angle = 0.100586 pi
    12'b000011010000: begin  real1=16'b0011110011000101; imag1=16'b0001010000010011;  end  // angle = 0.101563 pi
    12'b000011010010: begin  real1=16'b0011110010110101; imag1=16'b0001010001000011;  end  // angle = 0.102539 pi
    12'b000011010100: begin  real1=16'b0011110010100101; imag1=16'b0001010001110011;  end  // angle = 0.103516 pi
    12'b000011010110: begin  real1=16'b0011110010010101; imag1=16'b0001010010100010;  end  // angle = 0.104492 pi
    12'b000011011000: begin  real1=16'b0011110010000101; imag1=16'b0001010011010010;  end  // angle = 0.105469 pi
    12'b000011011010: begin  real1=16'b0011110001110100; imag1=16'b0001010100000001;  end  // angle = 0.106445 pi
    12'b000011011100: begin  real1=16'b0011110001100100; imag1=16'b0001010100110001;  end  // angle = 0.107422 pi
    12'b000011011110: begin  real1=16'b0011110001010011; imag1=16'b0001010101100000;  end  // angle = 0.108398 pi
    12'b000011100000: begin  real1=16'b0011110001000010; imag1=16'b0001010110010000;  end  // angle = 0.109375 pi
    12'b000011100010: begin  real1=16'b0011110000110001; imag1=16'b0001010110111111;  end  // angle = 0.110352 pi
    12'b000011100100: begin  real1=16'b0011110000100000; imag1=16'b0001010111101110;  end  // angle = 0.111328 pi
    12'b000011100110: begin  real1=16'b0011110000001111; imag1=16'b0001011000011101;  end  // angle = 0.112305 pi
    12'b000011101000: begin  real1=16'b0011101111111101; imag1=16'b0001011001001100;  end  // angle = 0.113281 pi
    12'b000011101010: begin  real1=16'b0011101111101100; imag1=16'b0001011001111100;  end  // angle = 0.114258 pi
    12'b000011101100: begin  real1=16'b0011101111011010; imag1=16'b0001011010101011;  end  // angle = 0.115234 pi
    12'b000011101110: begin  real1=16'b0011101111001000; imag1=16'b0001011011011010;  end  // angle = 0.116211 pi
    12'b000011110000: begin  real1=16'b0011101110110110; imag1=16'b0001011100001001;  end  // angle = 0.117187 pi
    12'b000011110010: begin  real1=16'b0011101110100100; imag1=16'b0001011100110111;  end  // angle = 0.118164 pi
    12'b000011110100: begin  real1=16'b0011101110010010; imag1=16'b0001011101100110;  end  // angle = 0.119141 pi
    12'b000011110110: begin  real1=16'b0011101101111111; imag1=16'b0001011110010101;  end  // angle = 0.120117 pi
    12'b000011111000: begin  real1=16'b0011101101101101; imag1=16'b0001011111000100;  end  // angle = 0.121094 pi
    12'b000011111010: begin  real1=16'b0011101101011010; imag1=16'b0001011111110010;  end  // angle = 0.122070 pi
    12'b000011111100: begin  real1=16'b0011101101000111; imag1=16'b0001100000100001;  end  // angle = 0.123047 pi
    12'b000011111110: begin  real1=16'b0011101100110100; imag1=16'b0001100001001111;  end  // angle = 0.124023 pi
    12'b000100000000: begin  real1=16'b0011101100100001; imag1=16'b0001100001111110;  end  // angle = 0.125000 pi
    12'b000100000010: begin  real1=16'b0011101100001110; imag1=16'b0001100010101100;  end  // angle = 0.125977 pi
    12'b000100000100: begin  real1=16'b0011101011111010; imag1=16'b0001100011011011;  end  // angle = 0.126953 pi
    12'b000100000110: begin  real1=16'b0011101011100110; imag1=16'b0001100100001001;  end  // angle = 0.127930 pi
    12'b000100001000: begin  real1=16'b0011101011010011; imag1=16'b0001100100110111;  end  // angle = 0.128906 pi
    12'b000100001010: begin  real1=16'b0011101010111111; imag1=16'b0001100101100101;  end  // angle = 0.129883 pi
    12'b000100001100: begin  real1=16'b0011101010101011; imag1=16'b0001100110010011;  end  // angle = 0.130859 pi
    12'b000100001110: begin  real1=16'b0011101010010111; imag1=16'b0001100111000001;  end  // angle = 0.131836 pi
    12'b000100010000: begin  real1=16'b0011101010000010; imag1=16'b0001100111101111;  end  // angle = 0.132812 pi
    12'b000100010010: begin  real1=16'b0011101001101110; imag1=16'b0001101000011101;  end  // angle = 0.133789 pi
    12'b000100010100: begin  real1=16'b0011101001011001; imag1=16'b0001101001001011;  end  // angle = 0.134766 pi
    12'b000100010110: begin  real1=16'b0011101001000101; imag1=16'b0001101001111001;  end  // angle = 0.135742 pi
    12'b000100011000: begin  real1=16'b0011101000110000; imag1=16'b0001101010100111;  end  // angle = 0.136719 pi
    12'b000100011010: begin  real1=16'b0011101000011011; imag1=16'b0001101011010100;  end  // angle = 0.137695 pi
    12'b000100011100: begin  real1=16'b0011101000000110; imag1=16'b0001101100000010;  end  // angle = 0.138672 pi
    12'b000100011110: begin  real1=16'b0011100111110000; imag1=16'b0001101100110000;  end  // angle = 0.139648 pi
    12'b000100100000: begin  real1=16'b0011100111011011; imag1=16'b0001101101011101;  end  // angle = 0.140625 pi
    12'b000100100010: begin  real1=16'b0011100111000101; imag1=16'b0001101110001010;  end  // angle = 0.141602 pi
    12'b000100100100: begin  real1=16'b0011100110110000; imag1=16'b0001101110111000;  end  // angle = 0.142578 pi
    12'b000100100110: begin  real1=16'b0011100110011010; imag1=16'b0001101111100101;  end  // angle = 0.143555 pi
    12'b000100101000: begin  real1=16'b0011100110000100; imag1=16'b0001110000010010;  end  // angle = 0.144531 pi
    12'b000100101010: begin  real1=16'b0011100101101110; imag1=16'b0001110000111111;  end  // angle = 0.145508 pi
    12'b000100101100: begin  real1=16'b0011100101011000; imag1=16'b0001110001101100;  end  // angle = 0.146484 pi
    12'b000100101110: begin  real1=16'b0011100101000001; imag1=16'b0001110010011001;  end  // angle = 0.147461 pi
    12'b000100110000: begin  real1=16'b0011100100101011; imag1=16'b0001110011000110;  end  // angle = 0.148438 pi
    12'b000100110010: begin  real1=16'b0011100100010100; imag1=16'b0001110011110011;  end  // angle = 0.149414 pi
    12'b000100110100: begin  real1=16'b0011100011111101; imag1=16'b0001110100100000;  end  // angle = 0.150391 pi
    12'b000100110110: begin  real1=16'b0011100011100110; imag1=16'b0001110101001101;  end  // angle = 0.151367 pi
    12'b000100111000: begin  real1=16'b0011100011001111; imag1=16'b0001110101111001;  end  // angle = 0.152344 pi
    12'b000100111010: begin  real1=16'b0011100010111000; imag1=16'b0001110110100110;  end  // angle = 0.153320 pi
    12'b000100111100: begin  real1=16'b0011100010100001; imag1=16'b0001110111010011;  end  // angle = 0.154297 pi
    12'b000100111110: begin  real1=16'b0011100010001001; imag1=16'b0001110111111111;  end  // angle = 0.155273 pi
    12'b000101000000: begin  real1=16'b0011100001110001; imag1=16'b0001111000101011;  end  // angle = 0.156250 pi
    12'b000101000010: begin  real1=16'b0011100001011010; imag1=16'b0001111001011000;  end  // angle = 0.157227 pi
    12'b000101000100: begin  real1=16'b0011100001000010; imag1=16'b0001111010000100;  end  // angle = 0.158203 pi
    12'b000101000110: begin  real1=16'b0011100000101010; imag1=16'b0001111010110000;  end  // angle = 0.159180 pi
    12'b000101001000: begin  real1=16'b0011100000010010; imag1=16'b0001111011011100;  end  // angle = 0.160156 pi
    12'b000101001010: begin  real1=16'b0011011111111001; imag1=16'b0001111100001000;  end  // angle = 0.161133 pi
    12'b000101001100: begin  real1=16'b0011011111100001; imag1=16'b0001111100110100;  end  // angle = 0.162109 pi
    12'b000101001110: begin  real1=16'b0011011111001000; imag1=16'b0001111101100000;  end  // angle = 0.163086 pi
    12'b000101010000: begin  real1=16'b0011011110110000; imag1=16'b0001111110001100;  end  // angle = 0.164062 pi
    12'b000101010010: begin  real1=16'b0011011110010111; imag1=16'b0001111110110111;  end  // angle = 0.165039 pi
    12'b000101010100: begin  real1=16'b0011011101111110; imag1=16'b0001111111100011;  end  // angle = 0.166016 pi
    12'b000101010110: begin  real1=16'b0011011101100101; imag1=16'b0010000000001111;  end  // angle = 0.166992 pi
    12'b000101011000: begin  real1=16'b0011011101001011; imag1=16'b0010000000111010;  end  // angle = 0.167969 pi
    12'b000101011010: begin  real1=16'b0011011100110010; imag1=16'b0010000001100101;  end  // angle = 0.168945 pi
    12'b000101011100: begin  real1=16'b0011011100011000; imag1=16'b0010000010010001;  end  // angle = 0.169922 pi
    12'b000101011110: begin  real1=16'b0011011011111111; imag1=16'b0010000010111100;  end  // angle = 0.170898 pi
    12'b000101100000: begin  real1=16'b0011011011100101; imag1=16'b0010000011100111;  end  // angle = 0.171875 pi
    12'b000101100010: begin  real1=16'b0011011011001011; imag1=16'b0010000100010010;  end  // angle = 0.172852 pi
    12'b000101100100: begin  real1=16'b0011011010110001; imag1=16'b0010000100111101;  end  // angle = 0.173828 pi
    12'b000101100110: begin  real1=16'b0011011010010111; imag1=16'b0010000101101000;  end  // angle = 0.174805 pi
    12'b000101101000: begin  real1=16'b0011011001111101; imag1=16'b0010000110010011;  end  // angle = 0.175781 pi
    12'b000101101010: begin  real1=16'b0011011001100010; imag1=16'b0010000110111110;  end  // angle = 0.176758 pi
    12'b000101101100: begin  real1=16'b0011011001001000; imag1=16'b0010000111101000;  end  // angle = 0.177734 pi
    12'b000101101110: begin  real1=16'b0011011000101101; imag1=16'b0010001000010011;  end  // angle = 0.178711 pi
    12'b000101110000: begin  real1=16'b0011011000010010; imag1=16'b0010001000111101;  end  // angle = 0.179688 pi
    12'b000101110010: begin  real1=16'b0011010111110111; imag1=16'b0010001001101000;  end  // angle = 0.180664 pi
    12'b000101110100: begin  real1=16'b0011010111011100; imag1=16'b0010001010010010;  end  // angle = 0.181641 pi
    12'b000101110110: begin  real1=16'b0011010111000001; imag1=16'b0010001010111100;  end  // angle = 0.182617 pi
    12'b000101111000: begin  real1=16'b0011010110100101; imag1=16'b0010001011100111;  end  // angle = 0.183594 pi
    12'b000101111010: begin  real1=16'b0011010110001010; imag1=16'b0010001100010001;  end  // angle = 0.184570 pi
    12'b000101111100: begin  real1=16'b0011010101101110; imag1=16'b0010001100111011;  end  // angle = 0.185547 pi
    12'b000101111110: begin  real1=16'b0011010101010011; imag1=16'b0010001101100101;  end  // angle = 0.186523 pi
    12'b000110000000: begin  real1=16'b0011010100110111; imag1=16'b0010001110001110;  end  // angle = 0.187500 pi
    12'b000110000010: begin  real1=16'b0011010100011011; imag1=16'b0010001110111000;  end  // angle = 0.188477 pi
    12'b000110000100: begin  real1=16'b0011010011111111; imag1=16'b0010001111100010;  end  // angle = 0.189453 pi
    12'b000110000110: begin  real1=16'b0011010011100010; imag1=16'b0010010000001011;  end  // angle = 0.190430 pi
    12'b000110001000: begin  real1=16'b0011010011000110; imag1=16'b0010010000110101;  end  // angle = 0.191406 pi
    12'b000110001010: begin  real1=16'b0011010010101010; imag1=16'b0010010001011110;  end  // angle = 0.192383 pi
    12'b000110001100: begin  real1=16'b0011010010001101; imag1=16'b0010010010001000;  end  // angle = 0.193359 pi
    12'b000110001110: begin  real1=16'b0011010001110000; imag1=16'b0010010010110001;  end  // angle = 0.194336 pi
    12'b000110010000: begin  real1=16'b0011010001010011; imag1=16'b0010010011011010;  end  // angle = 0.195312 pi
    12'b000110010010: begin  real1=16'b0011010000110110; imag1=16'b0010010100000011;  end  // angle = 0.196289 pi
    12'b000110010100: begin  real1=16'b0011010000011001; imag1=16'b0010010100101100;  end  // angle = 0.197266 pi
    12'b000110010110: begin  real1=16'b0011001111111100; imag1=16'b0010010101010101;  end  // angle = 0.198242 pi
    12'b000110011000: begin  real1=16'b0011001111011111; imag1=16'b0010010101111110;  end  // angle = 0.199219 pi
    12'b000110011010: begin  real1=16'b0011001111000001; imag1=16'b0010010110100110;  end  // angle = 0.200195 pi
    12'b000110011100: begin  real1=16'b0011001110100011; imag1=16'b0010010111001111;  end  // angle = 0.201172 pi
    12'b000110011110: begin  real1=16'b0011001110000110; imag1=16'b0010010111111000;  end  // angle = 0.202148 pi
    12'b000110100000: begin  real1=16'b0011001101101000; imag1=16'b0010011000100000;  end  // angle = 0.203125 pi
    12'b000110100010: begin  real1=16'b0011001101001010; imag1=16'b0010011001001000;  end  // angle = 0.204102 pi
    12'b000110100100: begin  real1=16'b0011001100101100; imag1=16'b0010011001110001;  end  // angle = 0.205078 pi
    12'b000110100110: begin  real1=16'b0011001100001101; imag1=16'b0010011010011001;  end  // angle = 0.206055 pi
    12'b000110101000: begin  real1=16'b0011001011101111; imag1=16'b0010011011000001;  end  // angle = 0.207031 pi
    12'b000110101010: begin  real1=16'b0011001011010000; imag1=16'b0010011011101001;  end  // angle = 0.208008 pi
    12'b000110101100: begin  real1=16'b0011001010110010; imag1=16'b0010011100010001;  end  // angle = 0.208984 pi
    12'b000110101110: begin  real1=16'b0011001010010011; imag1=16'b0010011100111000;  end  // angle = 0.209961 pi
    12'b000110110000: begin  real1=16'b0011001001110100; imag1=16'b0010011101100000;  end  // angle = 0.210938 pi
    12'b000110110010: begin  real1=16'b0011001001010101; imag1=16'b0010011110001000;  end  // angle = 0.211914 pi
    12'b000110110100: begin  real1=16'b0011001000110110; imag1=16'b0010011110101111;  end  // angle = 0.212891 pi
    12'b000110110110: begin  real1=16'b0011001000010111; imag1=16'b0010011111010110;  end  // angle = 0.213867 pi
    12'b000110111000: begin  real1=16'b0011000111111000; imag1=16'b0010011111111110;  end  // angle = 0.214844 pi
    12'b000110111010: begin  real1=16'b0011000111011000; imag1=16'b0010100000100101;  end  // angle = 0.215820 pi
    12'b000110111100: begin  real1=16'b0011000110111001; imag1=16'b0010100001001100;  end  // angle = 0.216797 pi
    12'b000110111110: begin  real1=16'b0011000110011001; imag1=16'b0010100001110011;  end  // angle = 0.217773 pi
    12'b000111000000: begin  real1=16'b0011000101111001; imag1=16'b0010100010011010;  end  // angle = 0.218750 pi
    12'b000111000010: begin  real1=16'b0011000101011001; imag1=16'b0010100011000001;  end  // angle = 0.219727 pi
    12'b000111000100: begin  real1=16'b0011000100111001; imag1=16'b0010100011100111;  end  // angle = 0.220703 pi
    12'b000111000110: begin  real1=16'b0011000100011001; imag1=16'b0010100100001110;  end  // angle = 0.221680 pi
    12'b000111001000: begin  real1=16'b0011000011111001; imag1=16'b0010100100110101;  end  // angle = 0.222656 pi
    12'b000111001010: begin  real1=16'b0011000011011000; imag1=16'b0010100101011011;  end  // angle = 0.223633 pi
    12'b000111001100: begin  real1=16'b0011000010111000; imag1=16'b0010100110000001;  end  // angle = 0.224609 pi
    12'b000111001110: begin  real1=16'b0011000010010111; imag1=16'b0010100110100111;  end  // angle = 0.225586 pi
    12'b000111010000: begin  real1=16'b0011000001110110; imag1=16'b0010100111001110;  end  // angle = 0.226562 pi
    12'b000111010010: begin  real1=16'b0011000001010101; imag1=16'b0010100111110100;  end  // angle = 0.227539 pi
    12'b000111010100: begin  real1=16'b0011000000110100; imag1=16'b0010101000011010;  end  // angle = 0.228516 pi
    12'b000111010110: begin  real1=16'b0011000000010011; imag1=16'b0010101000111111;  end  // angle = 0.229492 pi
    12'b000111011000: begin  real1=16'b0010111111110010; imag1=16'b0010101001100101;  end  // angle = 0.230469 pi
    12'b000111011010: begin  real1=16'b0010111111010000; imag1=16'b0010101010001011;  end  // angle = 0.231445 pi
    12'b000111011100: begin  real1=16'b0010111110101111; imag1=16'b0010101010110000;  end  // angle = 0.232422 pi
    12'b000111011110: begin  real1=16'b0010111110001101; imag1=16'b0010101011010110;  end  // angle = 0.233398 pi
    12'b000111100000: begin  real1=16'b0010111101101100; imag1=16'b0010101011111011;  end  // angle = 0.234375 pi
    12'b000111100010: begin  real1=16'b0010111101001010; imag1=16'b0010101100100000;  end  // angle = 0.235352 pi
    12'b000111100100: begin  real1=16'b0010111100101000; imag1=16'b0010101101000101;  end  // angle = 0.236328 pi
    12'b000111100110: begin  real1=16'b0010111100000110; imag1=16'b0010101101101010;  end  // angle = 0.237305 pi
    12'b000111101000: begin  real1=16'b0010111011100100; imag1=16'b0010101110001111;  end  // angle = 0.238281 pi
    12'b000111101010: begin  real1=16'b0010111011000010; imag1=16'b0010101110110100;  end  // angle = 0.239258 pi
    12'b000111101100: begin  real1=16'b0010111010011111; imag1=16'b0010101111011000;  end  // angle = 0.240234 pi
    12'b000111101110: begin  real1=16'b0010111001111101; imag1=16'b0010101111111101;  end  // angle = 0.241211 pi
    12'b000111110000: begin  real1=16'b0010111001011010; imag1=16'b0010110000100001;  end  // angle = 0.242188 pi
    12'b000111110010: begin  real1=16'b0010111000110111; imag1=16'b0010110001000110;  end  // angle = 0.243164 pi
    12'b000111110100: begin  real1=16'b0010111000010101; imag1=16'b0010110001101010;  end  // angle = 0.244141 pi
    12'b000111110110: begin  real1=16'b0010110111110010; imag1=16'b0010110010001110;  end  // angle = 0.245117 pi
    12'b000111111000: begin  real1=16'b0010110111001111; imag1=16'b0010110010110010;  end  // angle = 0.246094 pi
    12'b000111111010: begin  real1=16'b0010110110101011; imag1=16'b0010110011010110;  end  // angle = 0.247070 pi
    12'b000111111100: begin  real1=16'b0010110110001000; imag1=16'b0010110011111010;  end  // angle = 0.248047 pi
    12'b000111111110: begin  real1=16'b0010110101100101; imag1=16'b0010110100011110;  end  // angle = 0.249023 pi
    12'b001000000000: begin  real1=16'b0010110101000001; imag1=16'b0010110101000001;  end  // angle = 0.250000 pi
endcase
end


endmodule
