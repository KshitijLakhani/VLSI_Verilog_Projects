module ComplexExponential (
input [11:0] in_theta,
output reg [15:0] out_real,
output reg [15:0] out_imag);

always @(in_theta) begin
 case (in_theta)
 12'b000000000000: begin out_real=16'b0100000000000000; out_imag=16'b0000000000000000; end // in_theta = 0.000000 pi
 12'b000000000001: begin out_real=16'b0100000000000000; out_imag=16'b0000000000011001; end // in_theta = 0.000488 pi
 12'b000000000010: begin out_real=16'b0100000000000000; out_imag=16'b0000000000110010; end // in_theta = 0.000977 pi
 12'b000000000011: begin out_real=16'b0100000000000000; out_imag=16'b0000000001001011; end // in_theta = 0.001465 pi
 12'b000000000100: begin out_real=16'b0100000000000000; out_imag=16'b0000000001100101; end // in_theta = 0.001953 pi
 12'b000000000101: begin out_real=16'b0100000000000000; out_imag=16'b0000000001111110; end // in_theta = 0.002441 pi
 12'b000000000110: begin out_real=16'b0011111111111111; out_imag=16'b0000000010010111; end // in_theta = 0.002930 pi
 12'b000000000111: begin out_real=16'b0011111111111111; out_imag=16'b0000000010110000; end // in_theta = 0.003418 pi
 12'b000000001000: begin out_real=16'b0011111111111111; out_imag=16'b0000000011001001; end // in_theta = 0.003906 pi
 12'b000000001001: begin out_real=16'b0011111111111110; out_imag=16'b0000000011100010; end // in_theta = 0.004395 pi
 12'b000000001010: begin out_real=16'b0011111111111110; out_imag=16'b0000000011111011; end // in_theta = 0.004883 pi
 12'b000000001011: begin out_real=16'b0011111111111110; out_imag=16'b0000000100010100; end // in_theta = 0.005371 pi
 12'b000000001100: begin out_real=16'b0011111111111101; out_imag=16'b0000000100101110; end // in_theta = 0.005859 pi
 12'b000000001101: begin out_real=16'b0011111111111101; out_imag=16'b0000000101000111; end // in_theta = 0.006348 pi
 12'b000000001110: begin out_real=16'b0011111111111100; out_imag=16'b0000000101100000; end // in_theta = 0.006836 pi
 12'b000000001111: begin out_real=16'b0011111111111100; out_imag=16'b0000000101111001; end // in_theta = 0.007324 pi
 12'b000000010000: begin out_real=16'b0011111111111011; out_imag=16'b0000000110010010; end // in_theta = 0.007813 pi
 12'b000000010001: begin out_real=16'b0011111111111010; out_imag=16'b0000000110101011; end // in_theta = 0.008301 pi
 12'b000000010010: begin out_real=16'b0011111111111010; out_imag=16'b0000000111000100; end // in_theta = 0.008789 pi
 12'b000000010011: begin out_real=16'b0011111111111001; out_imag=16'b0000000111011101; end // in_theta = 0.009277 pi
 12'b000000010100: begin out_real=16'b0011111111111000; out_imag=16'b0000000111110111; end // in_theta = 0.009766 pi
 12'b000000010101: begin out_real=16'b0011111111110111; out_imag=16'b0000001000010000; end // in_theta = 0.010254 pi
 12'b000000010110: begin out_real=16'b0011111111110111; out_imag=16'b0000001000101001; end // in_theta = 0.010742 pi
 12'b000000010111: begin out_real=16'b0011111111110110; out_imag=16'b0000001001000010; end // in_theta = 0.011230 pi
 12'b000000011000: begin out_real=16'b0011111111110101; out_imag=16'b0000001001011011; end // in_theta = 0.011719 pi
 12'b000000011001: begin out_real=16'b0011111111110100; out_imag=16'b0000001001110100; end // in_theta = 0.012207 pi
 12'b000000011010: begin out_real=16'b0011111111110011; out_imag=16'b0000001010001101; end // in_theta = 0.012695 pi
 12'b000000011011: begin out_real=16'b0011111111110010; out_imag=16'b0000001010100110; end // in_theta = 0.013184 pi
 12'b000000011100: begin out_real=16'b0011111111110001; out_imag=16'b0000001011000000; end // in_theta = 0.013672 pi
 12'b000000011101: begin out_real=16'b0011111111110000; out_imag=16'b0000001011011001; end // in_theta = 0.014160 pi
 12'b000000011110: begin out_real=16'b0011111111101111; out_imag=16'b0000001011110010; end // in_theta = 0.014648 pi
 12'b000000011111: begin out_real=16'b0011111111101101; out_imag=16'b0000001100001011; end // in_theta = 0.015137 pi
 12'b000000100000: begin out_real=16'b0011111111101100; out_imag=16'b0000001100100100; end // in_theta = 0.015625 pi
 12'b000000100001: begin out_real=16'b0011111111101011; out_imag=16'b0000001100111101; end // in_theta = 0.016113 pi
 12'b000000100010: begin out_real=16'b0011111111101010; out_imag=16'b0000001101010110; end // in_theta = 0.016602 pi
 12'b000000100011: begin out_real=16'b0011111111101000; out_imag=16'b0000001101101111; end // in_theta = 0.017090 pi
 12'b000000100100: begin out_real=16'b0011111111100111; out_imag=16'b0000001110001000; end // in_theta = 0.017578 pi
 12'b000000100101: begin out_real=16'b0011111111100110; out_imag=16'b0000001110100001; end // in_theta = 0.018066 pi
 12'b000000100110: begin out_real=16'b0011111111100100; out_imag=16'b0000001110111011; end // in_theta = 0.018555 pi
 12'b000000100111: begin out_real=16'b0011111111100011; out_imag=16'b0000001111010100; end // in_theta = 0.019043 pi
 12'b000000101000: begin out_real=16'b0011111111100001; out_imag=16'b0000001111101101; end // in_theta = 0.019531 pi
 12'b000000101001: begin out_real=16'b0011111111100000; out_imag=16'b0000010000000110; end // in_theta = 0.020020 pi
 12'b000000101010: begin out_real=16'b0011111111011110; out_imag=16'b0000010000011111; end // in_theta = 0.020508 pi
 12'b000000101011: begin out_real=16'b0011111111011100; out_imag=16'b0000010000111000; end // in_theta = 0.020996 pi
 12'b000000101100: begin out_real=16'b0011111111011011; out_imag=16'b0000010001010001; end // in_theta = 0.021484 pi
 12'b000000101101: begin out_real=16'b0011111111011001; out_imag=16'b0000010001101010; end // in_theta = 0.021973 pi
 12'b000000101110: begin out_real=16'b0011111111010111; out_imag=16'b0000010010000011; end // in_theta = 0.022461 pi
 12'b000000101111: begin out_real=16'b0011111111010101; out_imag=16'b0000010010011100; end // in_theta = 0.022949 pi
 12'b000000110000: begin out_real=16'b0011111111010100; out_imag=16'b0000010010110101; end // in_theta = 0.023438 pi
 12'b000000110001: begin out_real=16'b0011111111010010; out_imag=16'b0000010011001110; end // in_theta = 0.023926 pi
 12'b000000110010: begin out_real=16'b0011111111010000; out_imag=16'b0000010011100111; end // in_theta = 0.024414 pi
 12'b000000110011: begin out_real=16'b0011111111001110; out_imag=16'b0000010100000000; end // in_theta = 0.024902 pi
 12'b000000110100: begin out_real=16'b0011111111001100; out_imag=16'b0000010100011010; end // in_theta = 0.025391 pi
 12'b000000110101: begin out_real=16'b0011111111001010; out_imag=16'b0000010100110011; end // in_theta = 0.025879 pi
 12'b000000110110: begin out_real=16'b0011111111001000; out_imag=16'b0000010101001100; end // in_theta = 0.026367 pi
 12'b000000110111: begin out_real=16'b0011111111000110; out_imag=16'b0000010101100101; end // in_theta = 0.026855 pi
 12'b000000111000: begin out_real=16'b0011111111000100; out_imag=16'b0000010101111110; end // in_theta = 0.027344 pi
 12'b000000111001: begin out_real=16'b0011111111000001; out_imag=16'b0000010110010111; end // in_theta = 0.027832 pi
 12'b000000111010: begin out_real=16'b0011111110111111; out_imag=16'b0000010110110000; end // in_theta = 0.028320 pi
 12'b000000111011: begin out_real=16'b0011111110111101; out_imag=16'b0000010111001001; end // in_theta = 0.028809 pi
 12'b000000111100: begin out_real=16'b0011111110111011; out_imag=16'b0000010111100010; end // in_theta = 0.029297 pi
 12'b000000111101: begin out_real=16'b0011111110111000; out_imag=16'b0000010111111011; end // in_theta = 0.029785 pi
 12'b000000111110: begin out_real=16'b0011111110110110; out_imag=16'b0000011000010100; end // in_theta = 0.030273 pi
 12'b000000111111: begin out_real=16'b0011111110110100; out_imag=16'b0000011000101101; end // in_theta = 0.030762 pi
 12'b000001000000: begin out_real=16'b0011111110110001; out_imag=16'b0000011001000110; end // in_theta = 0.031250 pi
 12'b000001000001: begin out_real=16'b0011111110101111; out_imag=16'b0000011001011111; end // in_theta = 0.031738 pi
 12'b000001000010: begin out_real=16'b0011111110101100; out_imag=16'b0000011001111000; end // in_theta = 0.032227 pi
 12'b000001000011: begin out_real=16'b0011111110101010; out_imag=16'b0000011010010001; end // in_theta = 0.032715 pi
 12'b000001000100: begin out_real=16'b0011111110100111; out_imag=16'b0000011010101010; end // in_theta = 0.033203 pi
 12'b000001000101: begin out_real=16'b0011111110100100; out_imag=16'b0000011011000011; end // in_theta = 0.033691 pi
 12'b000001000110: begin out_real=16'b0011111110100010; out_imag=16'b0000011011011100; end // in_theta = 0.034180 pi
 12'b000001000111: begin out_real=16'b0011111110011111; out_imag=16'b0000011011110101; end // in_theta = 0.034668 pi
 12'b000001001000: begin out_real=16'b0011111110011100; out_imag=16'b0000011100001110; end // in_theta = 0.035156 pi
 12'b000001001001: begin out_real=16'b0011111110011001; out_imag=16'b0000011100100111; end // in_theta = 0.035645 pi
 12'b000001001010: begin out_real=16'b0011111110010111; out_imag=16'b0000011101000000; end // in_theta = 0.036133 pi
 12'b000001001011: begin out_real=16'b0011111110010100; out_imag=16'b0000011101011001; end // in_theta = 0.036621 pi
 12'b000001001100: begin out_real=16'b0011111110010001; out_imag=16'b0000011101110010; end // in_theta = 0.037109 pi
 12'b000001001101: begin out_real=16'b0011111110001110; out_imag=16'b0000011110001011; end // in_theta = 0.037598 pi
 12'b000001001110: begin out_real=16'b0011111110001011; out_imag=16'b0000011110100100; end // in_theta = 0.038086 pi
 12'b000001001111: begin out_real=16'b0011111110001000; out_imag=16'b0000011110111101; end // in_theta = 0.038574 pi
 12'b000001010000: begin out_real=16'b0011111110000101; out_imag=16'b0000011111010110; end // in_theta = 0.039063 pi
 12'b000001010001: begin out_real=16'b0011111110000010; out_imag=16'b0000011111101111; end // in_theta = 0.039551 pi
 12'b000001010010: begin out_real=16'b0011111101111111; out_imag=16'b0000100000000111; end // in_theta = 0.040039 pi
 12'b000001010011: begin out_real=16'b0011111101111011; out_imag=16'b0000100000100000; end // in_theta = 0.040527 pi
 12'b000001010100: begin out_real=16'b0011111101111000; out_imag=16'b0000100000111001; end // in_theta = 0.041016 pi
 12'b000001010101: begin out_real=16'b0011111101110101; out_imag=16'b0000100001010010; end // in_theta = 0.041504 pi
 12'b000001010110: begin out_real=16'b0011111101110010; out_imag=16'b0000100001101011; end // in_theta = 0.041992 pi
 12'b000001010111: begin out_real=16'b0011111101101110; out_imag=16'b0000100010000100; end // in_theta = 0.042480 pi
 12'b000001011000: begin out_real=16'b0011111101101011; out_imag=16'b0000100010011101; end // in_theta = 0.042969 pi
 12'b000001011001: begin out_real=16'b0011111101101000; out_imag=16'b0000100010110110; end // in_theta = 0.043457 pi
 12'b000001011010: begin out_real=16'b0011111101100100; out_imag=16'b0000100011001111; end // in_theta = 0.043945 pi
 12'b000001011011: begin out_real=16'b0011111101100001; out_imag=16'b0000100011101000; end // in_theta = 0.044434 pi
 12'b000001011100: begin out_real=16'b0011111101011101; out_imag=16'b0000100100000001; end // in_theta = 0.044922 pi
 12'b000001011101: begin out_real=16'b0011111101011010; out_imag=16'b0000100100011001; end // in_theta = 0.045410 pi
 12'b000001011110: begin out_real=16'b0011111101010110; out_imag=16'b0000100100110010; end // in_theta = 0.045898 pi
 12'b000001011111: begin out_real=16'b0011111101010010; out_imag=16'b0000100101001011; end // in_theta = 0.046387 pi
 12'b000001100000: begin out_real=16'b0011111101001111; out_imag=16'b0000100101100100; end // in_theta = 0.046875 pi
 12'b000001100001: begin out_real=16'b0011111101001011; out_imag=16'b0000100101111101; end // in_theta = 0.047363 pi
 12'b000001100010: begin out_real=16'b0011111101000111; out_imag=16'b0000100110010110; end // in_theta = 0.047852 pi
 12'b000001100011: begin out_real=16'b0011111101000011; out_imag=16'b0000100110101111; end // in_theta = 0.048340 pi
 12'b000001100100: begin out_real=16'b0011111101000000; out_imag=16'b0000100111000111; end // in_theta = 0.048828 pi
 12'b000001100101: begin out_real=16'b0011111100111100; out_imag=16'b0000100111100000; end // in_theta = 0.049316 pi
 12'b000001100110: begin out_real=16'b0011111100111000; out_imag=16'b0000100111111001; end // in_theta = 0.049805 pi
 12'b000001100111: begin out_real=16'b0011111100110100; out_imag=16'b0000101000010010; end // in_theta = 0.050293 pi
 12'b000001101000: begin out_real=16'b0011111100110000; out_imag=16'b0000101000101011; end // in_theta = 0.050781 pi
 12'b000001101001: begin out_real=16'b0011111100101100; out_imag=16'b0000101001000100; end // in_theta = 0.051270 pi
 12'b000001101010: begin out_real=16'b0011111100101000; out_imag=16'b0000101001011100; end // in_theta = 0.051758 pi
 12'b000001101011: begin out_real=16'b0011111100100100; out_imag=16'b0000101001110101; end // in_theta = 0.052246 pi
 12'b000001101100: begin out_real=16'b0011111100100000; out_imag=16'b0000101010001110; end // in_theta = 0.052734 pi
 12'b000001101101: begin out_real=16'b0011111100011100; out_imag=16'b0000101010100111; end // in_theta = 0.053223 pi
 12'b000001101110: begin out_real=16'b0011111100010111; out_imag=16'b0000101011000000; end // in_theta = 0.053711 pi
 12'b000001101111: begin out_real=16'b0011111100010011; out_imag=16'b0000101011011000; end // in_theta = 0.054199 pi
 12'b000001110000: begin out_real=16'b0011111100001111; out_imag=16'b0000101011110001; end // in_theta = 0.054688 pi
 12'b000001110001: begin out_real=16'b0011111100001010; out_imag=16'b0000101100001010; end // in_theta = 0.055176 pi
 12'b000001110010: begin out_real=16'b0011111100000110; out_imag=16'b0000101100100011; end // in_theta = 0.055664 pi
 12'b000001110011: begin out_real=16'b0011111100000010; out_imag=16'b0000101100111011; end // in_theta = 0.056152 pi
 12'b000001110100: begin out_real=16'b0011111011111101; out_imag=16'b0000101101010100; end // in_theta = 0.056641 pi
 12'b000001110101: begin out_real=16'b0011111011111001; out_imag=16'b0000101101101101; end // in_theta = 0.057129 pi
 12'b000001110110: begin out_real=16'b0011111011110100; out_imag=16'b0000101110000101; end // in_theta = 0.057617 pi
 12'b000001110111: begin out_real=16'b0011111011110000; out_imag=16'b0000101110011110; end // in_theta = 0.058105 pi
 12'b000001111000: begin out_real=16'b0011111011101011; out_imag=16'b0000101110110111; end // in_theta = 0.058594 pi
 12'b000001111001: begin out_real=16'b0011111011100111; out_imag=16'b0000101111010000; end // in_theta = 0.059082 pi
 12'b000001111010: begin out_real=16'b0011111011100010; out_imag=16'b0000101111101000; end // in_theta = 0.059570 pi
 12'b000001111011: begin out_real=16'b0011111011011101; out_imag=16'b0000110000000001; end // in_theta = 0.060059 pi
 12'b000001111100: begin out_real=16'b0011111011011000; out_imag=16'b0000110000011010; end // in_theta = 0.060547 pi
 12'b000001111101: begin out_real=16'b0011111011010100; out_imag=16'b0000110000110010; end // in_theta = 0.061035 pi
 12'b000001111110: begin out_real=16'b0011111011001111; out_imag=16'b0000110001001011; end // in_theta = 0.061523 pi
 12'b000001111111: begin out_real=16'b0011111011001010; out_imag=16'b0000110001100100; end // in_theta = 0.062012 pi
 12'b000010000000: begin out_real=16'b0011111011000101; out_imag=16'b0000110001111100; end // in_theta = 0.062500 pi
 12'b000010000001: begin out_real=16'b0011111011000000; out_imag=16'b0000110010010101; end // in_theta = 0.062988 pi
 12'b000010000010: begin out_real=16'b0011111010111011; out_imag=16'b0000110010101110; end // in_theta = 0.063477 pi
 12'b000010000011: begin out_real=16'b0011111010110110; out_imag=16'b0000110011000110; end // in_theta = 0.063965 pi
 12'b000010000100: begin out_real=16'b0011111010110001; out_imag=16'b0000110011011111; end // in_theta = 0.064453 pi
 12'b000010000101: begin out_real=16'b0011111010101100; out_imag=16'b0000110011111000; end // in_theta = 0.064941 pi
 12'b000010000110: begin out_real=16'b0011111010100111; out_imag=16'b0000110100010000; end // in_theta = 0.065430 pi
 12'b000010000111: begin out_real=16'b0011111010100010; out_imag=16'b0000110100101001; end // in_theta = 0.065918 pi
 12'b000010001000: begin out_real=16'b0011111010011101; out_imag=16'b0000110101000001; end // in_theta = 0.066406 pi
 12'b000010001001: begin out_real=16'b0011111010011000; out_imag=16'b0000110101011010; end // in_theta = 0.066895 pi
 12'b000010001010: begin out_real=16'b0011111010010010; out_imag=16'b0000110101110010; end // in_theta = 0.067383 pi
 12'b000010001011: begin out_real=16'b0011111010001101; out_imag=16'b0000110110001011; end // in_theta = 0.067871 pi
 12'b000010001100: begin out_real=16'b0011111010001000; out_imag=16'b0000110110100100; end // in_theta = 0.068359 pi
 12'b000010001101: begin out_real=16'b0011111010000010; out_imag=16'b0000110110111100; end // in_theta = 0.068848 pi
 12'b000010001110: begin out_real=16'b0011111001111101; out_imag=16'b0000110111010101; end // in_theta = 0.069336 pi
 12'b000010001111: begin out_real=16'b0011111001110111; out_imag=16'b0000110111101101; end // in_theta = 0.069824 pi
 12'b000010010000: begin out_real=16'b0011111001110010; out_imag=16'b0000111000000110; end // in_theta = 0.070313 pi
 12'b000010010001: begin out_real=16'b0011111001101100; out_imag=16'b0000111000011110; end // in_theta = 0.070801 pi
 12'b000010010010: begin out_real=16'b0011111001100111; out_imag=16'b0000111000110111; end // in_theta = 0.071289 pi
 12'b000010010011: begin out_real=16'b0011111001100001; out_imag=16'b0000111001001111; end // in_theta = 0.071777 pi
 12'b000010010100: begin out_real=16'b0011111001011100; out_imag=16'b0000111001101000; end // in_theta = 0.072266 pi
 12'b000010010101: begin out_real=16'b0011111001010110; out_imag=16'b0000111010000000; end // in_theta = 0.072754 pi
 12'b000010010110: begin out_real=16'b0011111001010000; out_imag=16'b0000111010011001; end // in_theta = 0.073242 pi
 12'b000010010111: begin out_real=16'b0011111001001010; out_imag=16'b0000111010110001; end // in_theta = 0.073730 pi
 12'b000010011000: begin out_real=16'b0011111001000101; out_imag=16'b0000111011001010; end // in_theta = 0.074219 pi
 12'b000010011001: begin out_real=16'b0011111000111111; out_imag=16'b0000111011100010; end // in_theta = 0.074707 pi
 12'b000010011010: begin out_real=16'b0011111000111001; out_imag=16'b0000111011111011; end // in_theta = 0.075195 pi
 12'b000010011011: begin out_real=16'b0011111000110011; out_imag=16'b0000111100010011; end // in_theta = 0.075684 pi
 12'b000010011100: begin out_real=16'b0011111000101101; out_imag=16'b0000111100101011; end // in_theta = 0.076172 pi
 12'b000010011101: begin out_real=16'b0011111000100111; out_imag=16'b0000111101000100; end // in_theta = 0.076660 pi
 12'b000010011110: begin out_real=16'b0011111000100001; out_imag=16'b0000111101011100; end // in_theta = 0.077148 pi
 12'b000010011111: begin out_real=16'b0011111000011011; out_imag=16'b0000111101110101; end // in_theta = 0.077637 pi
 12'b000010100000: begin out_real=16'b0011111000010101; out_imag=16'b0000111110001101; end // in_theta = 0.078125 pi
 12'b000010100001: begin out_real=16'b0011111000001111; out_imag=16'b0000111110100101; end // in_theta = 0.078613 pi
 12'b000010100010: begin out_real=16'b0011111000001001; out_imag=16'b0000111110111110; end // in_theta = 0.079102 pi
 12'b000010100011: begin out_real=16'b0011111000000011; out_imag=16'b0000111111010110; end // in_theta = 0.079590 pi
 12'b000010100100: begin out_real=16'b0011110111111100; out_imag=16'b0000111111101110; end // in_theta = 0.080078 pi
 12'b000010100101: begin out_real=16'b0011110111110110; out_imag=16'b0001000000000111; end // in_theta = 0.080566 pi
 12'b000010100110: begin out_real=16'b0011110111110000; out_imag=16'b0001000000011111; end // in_theta = 0.081055 pi
 12'b000010100111: begin out_real=16'b0011110111101001; out_imag=16'b0001000000110111; end // in_theta = 0.081543 pi
 12'b000010101000: begin out_real=16'b0011110111100011; out_imag=16'b0001000001010000; end // in_theta = 0.082031 pi
 12'b000010101001: begin out_real=16'b0011110111011101; out_imag=16'b0001000001101000; end // in_theta = 0.082520 pi
 12'b000010101010: begin out_real=16'b0011110111010110; out_imag=16'b0001000010000000; end // in_theta = 0.083008 pi
 12'b000010101011: begin out_real=16'b0011110111010000; out_imag=16'b0001000010011001; end // in_theta = 0.083496 pi
 12'b000010101100: begin out_real=16'b0011110111001001; out_imag=16'b0001000010110001; end // in_theta = 0.083984 pi
 12'b000010101101: begin out_real=16'b0011110111000010; out_imag=16'b0001000011001001; end // in_theta = 0.084473 pi
 12'b000010101110: begin out_real=16'b0011110110111100; out_imag=16'b0001000011100001; end // in_theta = 0.084961 pi
 12'b000010101111: begin out_real=16'b0011110110110101; out_imag=16'b0001000011111010; end // in_theta = 0.085449 pi
 12'b000010110000: begin out_real=16'b0011110110101111; out_imag=16'b0001000100010010; end // in_theta = 0.085937 pi
 12'b000010110001: begin out_real=16'b0011110110101000; out_imag=16'b0001000100101010; end // in_theta = 0.086426 pi
 12'b000010110010: begin out_real=16'b0011110110100001; out_imag=16'b0001000101000010; end // in_theta = 0.086914 pi
 12'b000010110011: begin out_real=16'b0011110110011010; out_imag=16'b0001000101011010; end // in_theta = 0.087402 pi
 12'b000010110100: begin out_real=16'b0011110110010011; out_imag=16'b0001000101110011; end // in_theta = 0.087891 pi
 12'b000010110101: begin out_real=16'b0011110110001101; out_imag=16'b0001000110001011; end // in_theta = 0.088379 pi
 12'b000010110110: begin out_real=16'b0011110110000110; out_imag=16'b0001000110100011; end // in_theta = 0.088867 pi
 12'b000010110111: begin out_real=16'b0011110101111111; out_imag=16'b0001000110111011; end // in_theta = 0.089355 pi
 12'b000010111000: begin out_real=16'b0011110101111000; out_imag=16'b0001000111010011; end // in_theta = 0.089844 pi
 12'b000010111001: begin out_real=16'b0011110101110001; out_imag=16'b0001000111101011; end // in_theta = 0.090332 pi
 12'b000010111010: begin out_real=16'b0011110101101010; out_imag=16'b0001001000000100; end // in_theta = 0.090820 pi
 12'b000010111011: begin out_real=16'b0011110101100011; out_imag=16'b0001001000011100; end // in_theta = 0.091309 pi
 12'b000010111100: begin out_real=16'b0011110101011011; out_imag=16'b0001001000110100; end // in_theta = 0.091797 pi
 12'b000010111101: begin out_real=16'b0011110101010100; out_imag=16'b0001001001001100; end // in_theta = 0.092285 pi
 12'b000010111110: begin out_real=16'b0011110101001101; out_imag=16'b0001001001100100; end // in_theta = 0.092773 pi
 12'b000010111111: begin out_real=16'b0011110101000110; out_imag=16'b0001001001111100; end // in_theta = 0.093262 pi
 12'b000011000000: begin out_real=16'b0011110100111111; out_imag=16'b0001001010010100; end // in_theta = 0.093750 pi
 12'b000011000001: begin out_real=16'b0011110100110111; out_imag=16'b0001001010101100; end // in_theta = 0.094238 pi
 12'b000011000010: begin out_real=16'b0011110100110000; out_imag=16'b0001001011000100; end // in_theta = 0.094727 pi
 12'b000011000011: begin out_real=16'b0011110100101000; out_imag=16'b0001001011011100; end // in_theta = 0.095215 pi
 12'b000011000100: begin out_real=16'b0011110100100001; out_imag=16'b0001001011110100; end // in_theta = 0.095703 pi
 12'b000011000101: begin out_real=16'b0011110100011010; out_imag=16'b0001001100001100; end // in_theta = 0.096191 pi
 12'b000011000110: begin out_real=16'b0011110100010010; out_imag=16'b0001001100100100; end // in_theta = 0.096680 pi
 12'b000011000111: begin out_real=16'b0011110100001011; out_imag=16'b0001001100111100; end // in_theta = 0.097168 pi
 12'b000011001000: begin out_real=16'b0011110100000011; out_imag=16'b0001001101010100; end // in_theta = 0.097656 pi
 12'b000011001001: begin out_real=16'b0011110011111011; out_imag=16'b0001001101101100; end // in_theta = 0.098145 pi
 12'b000011001010: begin out_real=16'b0011110011110100; out_imag=16'b0001001110000100; end // in_theta = 0.098633 pi
 12'b000011001011: begin out_real=16'b0011110011101100; out_imag=16'b0001001110011100; end // in_theta = 0.099121 pi
 12'b000011001100: begin out_real=16'b0011110011100100; out_imag=16'b0001001110110100; end // in_theta = 0.099609 pi
 12'b000011001101: begin out_real=16'b0011110011011101; out_imag=16'b0001001111001100; end // in_theta = 0.100098 pi
 12'b000011001110: begin out_real=16'b0011110011010101; out_imag=16'b0001001111100100; end // in_theta = 0.100586 pi
 12'b000011001111: begin out_real=16'b0011110011001101; out_imag=16'b0001001111111011; end // in_theta = 0.101074 pi
 12'b000011010000: begin out_real=16'b0011110011000101; out_imag=16'b0001010000010011; end // in_theta = 0.101563 pi
 12'b000011010001: begin out_real=16'b0011110010111101; out_imag=16'b0001010000101011; end // in_theta = 0.102051 pi
 12'b000011010010: begin out_real=16'b0011110010110101; out_imag=16'b0001010001000011; end // in_theta = 0.102539 pi
 12'b000011010011: begin out_real=16'b0011110010101101; out_imag=16'b0001010001011011; end // in_theta = 0.103027 pi
 12'b000011010100: begin out_real=16'b0011110010100101; out_imag=16'b0001010001110011; end // in_theta = 0.103516 pi
 12'b000011010101: begin out_real=16'b0011110010011101; out_imag=16'b0001010010001011; end // in_theta = 0.104004 pi
 12'b000011010110: begin out_real=16'b0011110010010101; out_imag=16'b0001010010100010; end // in_theta = 0.104492 pi
 12'b000011010111: begin out_real=16'b0011110010001101; out_imag=16'b0001010010111010; end // in_theta = 0.104980 pi
 12'b000011011000: begin out_real=16'b0011110010000101; out_imag=16'b0001010011010010; end // in_theta = 0.105469 pi
 12'b000011011001: begin out_real=16'b0011110001111101; out_imag=16'b0001010011101010; end // in_theta = 0.105957 pi
 12'b000011011010: begin out_real=16'b0011110001110100; out_imag=16'b0001010100000001; end // in_theta = 0.106445 pi
 12'b000011011011: begin out_real=16'b0011110001101100; out_imag=16'b0001010100011001; end // in_theta = 0.106934 pi
 12'b000011011100: begin out_real=16'b0011110001100100; out_imag=16'b0001010100110001; end // in_theta = 0.107422 pi
 12'b000011011101: begin out_real=16'b0011110001011011; out_imag=16'b0001010101001001; end // in_theta = 0.107910 pi
 12'b000011011110: begin out_real=16'b0011110001010011; out_imag=16'b0001010101100000; end // in_theta = 0.108398 pi
 12'b000011011111: begin out_real=16'b0011110001001011; out_imag=16'b0001010101111000; end // in_theta = 0.108887 pi
 12'b000011100000: begin out_real=16'b0011110001000010; out_imag=16'b0001010110010000; end // in_theta = 0.109375 pi
 12'b000011100001: begin out_real=16'b0011110000111010; out_imag=16'b0001010110100111; end // in_theta = 0.109863 pi
 12'b000011100010: begin out_real=16'b0011110000110001; out_imag=16'b0001010110111111; end // in_theta = 0.110352 pi
 12'b000011100011: begin out_real=16'b0011110000101001; out_imag=16'b0001010111010111; end // in_theta = 0.110840 pi
 12'b000011100100: begin out_real=16'b0011110000100000; out_imag=16'b0001010111101110; end // in_theta = 0.111328 pi
 12'b000011100101: begin out_real=16'b0011110000010111; out_imag=16'b0001011000000110; end // in_theta = 0.111816 pi
 12'b000011100110: begin out_real=16'b0011110000001111; out_imag=16'b0001011000011101; end // in_theta = 0.112305 pi
 12'b000011100111: begin out_real=16'b0011110000000110; out_imag=16'b0001011000110101; end // in_theta = 0.112793 pi
 12'b000011101000: begin out_real=16'b0011101111111101; out_imag=16'b0001011001001100; end // in_theta = 0.113281 pi
 12'b000011101001: begin out_real=16'b0011101111110101; out_imag=16'b0001011001100100; end // in_theta = 0.113770 pi
 12'b000011101010: begin out_real=16'b0011101111101100; out_imag=16'b0001011001111100; end // in_theta = 0.114258 pi
 12'b000011101011: begin out_real=16'b0011101111100011; out_imag=16'b0001011010010011; end // in_theta = 0.114746 pi
 12'b000011101100: begin out_real=16'b0011101111011010; out_imag=16'b0001011010101011; end // in_theta = 0.115234 pi
 12'b000011101101: begin out_real=16'b0011101111010001; out_imag=16'b0001011011000010; end // in_theta = 0.115723 pi
 12'b000011101110: begin out_real=16'b0011101111001000; out_imag=16'b0001011011011010; end // in_theta = 0.116211 pi
 12'b000011101111: begin out_real=16'b0011101110111111; out_imag=16'b0001011011110001; end // in_theta = 0.116699 pi
 12'b000011110000: begin out_real=16'b0011101110110110; out_imag=16'b0001011100001001; end // in_theta = 0.117187 pi
 12'b000011110001: begin out_real=16'b0011101110101101; out_imag=16'b0001011100100000; end // in_theta = 0.117676 pi
 12'b000011110010: begin out_real=16'b0011101110100100; out_imag=16'b0001011100110111; end // in_theta = 0.118164 pi
 12'b000011110011: begin out_real=16'b0011101110011011; out_imag=16'b0001011101001111; end // in_theta = 0.118652 pi
 12'b000011110100: begin out_real=16'b0011101110010010; out_imag=16'b0001011101100110; end // in_theta = 0.119141 pi
 12'b000011110101: begin out_real=16'b0011101110001000; out_imag=16'b0001011101111110; end // in_theta = 0.119629 pi
 12'b000011110110: begin out_real=16'b0011101101111111; out_imag=16'b0001011110010101; end // in_theta = 0.120117 pi
 12'b000011110111: begin out_real=16'b0011101101110110; out_imag=16'b0001011110101100; end // in_theta = 0.120605 pi
 12'b000011111000: begin out_real=16'b0011101101101101; out_imag=16'b0001011111000100; end // in_theta = 0.121094 pi
 12'b000011111001: begin out_real=16'b0011101101100011; out_imag=16'b0001011111011011; end // in_theta = 0.121582 pi
 12'b000011111010: begin out_real=16'b0011101101011010; out_imag=16'b0001011111110010; end // in_theta = 0.122070 pi
 12'b000011111011: begin out_real=16'b0011101101010000; out_imag=16'b0001100000001010; end // in_theta = 0.122559 pi
 12'b000011111100: begin out_real=16'b0011101101000111; out_imag=16'b0001100000100001; end // in_theta = 0.123047 pi
 12'b000011111101: begin out_real=16'b0011101100111110; out_imag=16'b0001100000111000; end // in_theta = 0.123535 pi
 12'b000011111110: begin out_real=16'b0011101100110100; out_imag=16'b0001100001001111; end // in_theta = 0.124023 pi
 12'b000011111111: begin out_real=16'b0011101100101010; out_imag=16'b0001100001100111; end // in_theta = 0.124512 pi
 12'b000100000000: begin out_real=16'b0011101100100001; out_imag=16'b0001100001111110; end // in_theta = 0.125000 pi
 12'b000100000001: begin out_real=16'b0011101100010111; out_imag=16'b0001100010010101; end // in_theta = 0.125488 pi
 12'b000100000010: begin out_real=16'b0011101100001110; out_imag=16'b0001100010101100; end // in_theta = 0.125977 pi
 12'b000100000011: begin out_real=16'b0011101100000100; out_imag=16'b0001100011000011; end // in_theta = 0.126465 pi
 12'b000100000100: begin out_real=16'b0011101011111010; out_imag=16'b0001100011011011; end // in_theta = 0.126953 pi
 12'b000100000101: begin out_real=16'b0011101011110000; out_imag=16'b0001100011110010; end // in_theta = 0.127441 pi
 12'b000100000110: begin out_real=16'b0011101011100110; out_imag=16'b0001100100001001; end // in_theta = 0.127930 pi
 12'b000100000111: begin out_real=16'b0011101011011101; out_imag=16'b0001100100100000; end // in_theta = 0.128418 pi
 12'b000100001000: begin out_real=16'b0011101011010011; out_imag=16'b0001100100110111; end // in_theta = 0.128906 pi
 12'b000100001001: begin out_real=16'b0011101011001001; out_imag=16'b0001100101001110; end // in_theta = 0.129395 pi
 12'b000100001010: begin out_real=16'b0011101010111111; out_imag=16'b0001100101100101; end // in_theta = 0.129883 pi
 12'b000100001011: begin out_real=16'b0011101010110101; out_imag=16'b0001100101111100; end // in_theta = 0.130371 pi
 12'b000100001100: begin out_real=16'b0011101010101011; out_imag=16'b0001100110010011; end // in_theta = 0.130859 pi
 12'b000100001101: begin out_real=16'b0011101010100001; out_imag=16'b0001100110101010; end // in_theta = 0.131348 pi
 12'b000100001110: begin out_real=16'b0011101010010111; out_imag=16'b0001100111000001; end // in_theta = 0.131836 pi
 12'b000100001111: begin out_real=16'b0011101010001101; out_imag=16'b0001100111011000; end // in_theta = 0.132324 pi
 12'b000100010000: begin out_real=16'b0011101010000010; out_imag=16'b0001100111101111; end // in_theta = 0.132813 pi
 12'b000100010001: begin out_real=16'b0011101001111000; out_imag=16'b0001101000000110; end // in_theta = 0.133301 pi
 12'b000100010010: begin out_real=16'b0011101001101110; out_imag=16'b0001101000011101; end // in_theta = 0.133789 pi
 12'b000100010011: begin out_real=16'b0011101001100100; out_imag=16'b0001101000110100; end // in_theta = 0.134277 pi
 12'b000100010100: begin out_real=16'b0011101001011001; out_imag=16'b0001101001001011; end // in_theta = 0.134766 pi
 12'b000100010101: begin out_real=16'b0011101001001111; out_imag=16'b0001101001100010; end // in_theta = 0.135254 pi
 12'b000100010110: begin out_real=16'b0011101001000101; out_imag=16'b0001101001111001; end // in_theta = 0.135742 pi
 12'b000100010111: begin out_real=16'b0011101000111010; out_imag=16'b0001101010010000; end // in_theta = 0.136230 pi
 12'b000100011000: begin out_real=16'b0011101000110000; out_imag=16'b0001101010100111; end // in_theta = 0.136719 pi
 12'b000100011001: begin out_real=16'b0011101000100101; out_imag=16'b0001101010111110; end // in_theta = 0.137207 pi
 12'b000100011010: begin out_real=16'b0011101000011011; out_imag=16'b0001101011010100; end // in_theta = 0.137695 pi
 12'b000100011011: begin out_real=16'b0011101000010000; out_imag=16'b0001101011101011; end // in_theta = 0.138184 pi
 12'b000100011100: begin out_real=16'b0011101000000110; out_imag=16'b0001101100000010; end // in_theta = 0.138672 pi
 12'b000100011101: begin out_real=16'b0011100111111011; out_imag=16'b0001101100011001; end // in_theta = 0.139160 pi
 12'b000100011110: begin out_real=16'b0011100111110000; out_imag=16'b0001101100110000; end // in_theta = 0.139648 pi
 12'b000100011111: begin out_real=16'b0011100111100110; out_imag=16'b0001101101000110; end // in_theta = 0.140137 pi
 12'b000100100000: begin out_real=16'b0011100111011011; out_imag=16'b0001101101011101; end // in_theta = 0.140625 pi
 12'b000100100001: begin out_real=16'b0011100111010000; out_imag=16'b0001101101110100; end // in_theta = 0.141113 pi
 12'b000100100010: begin out_real=16'b0011100111000101; out_imag=16'b0001101110001010; end // in_theta = 0.141602 pi
 12'b000100100011: begin out_real=16'b0011100110111011; out_imag=16'b0001101110100001; end // in_theta = 0.142090 pi
 12'b000100100100: begin out_real=16'b0011100110110000; out_imag=16'b0001101110111000; end // in_theta = 0.142578 pi
 12'b000100100101: begin out_real=16'b0011100110100101; out_imag=16'b0001101111001110; end // in_theta = 0.143066 pi
 12'b000100100110: begin out_real=16'b0011100110011010; out_imag=16'b0001101111100101; end // in_theta = 0.143555 pi
 12'b000100100111: begin out_real=16'b0011100110001111; out_imag=16'b0001101111111100; end // in_theta = 0.144043 pi
 12'b000100101000: begin out_real=16'b0011100110000100; out_imag=16'b0001110000010010; end // in_theta = 0.144531 pi
 12'b000100101001: begin out_real=16'b0011100101111001; out_imag=16'b0001110000101001; end // in_theta = 0.145020 pi
 12'b000100101010: begin out_real=16'b0011100101101110; out_imag=16'b0001110000111111; end // in_theta = 0.145508 pi
 12'b000100101011: begin out_real=16'b0011100101100011; out_imag=16'b0001110001010110; end // in_theta = 0.145996 pi
 12'b000100101100: begin out_real=16'b0011100101011000; out_imag=16'b0001110001101100; end // in_theta = 0.146484 pi
 12'b000100101101: begin out_real=16'b0011100101001100; out_imag=16'b0001110010000011; end // in_theta = 0.146973 pi
 12'b000100101110: begin out_real=16'b0011100101000001; out_imag=16'b0001110010011001; end // in_theta = 0.147461 pi
 12'b000100101111: begin out_real=16'b0011100100110110; out_imag=16'b0001110010110000; end // in_theta = 0.147949 pi
 12'b000100110000: begin out_real=16'b0011100100101011; out_imag=16'b0001110011000110; end // in_theta = 0.148438 pi
 12'b000100110001: begin out_real=16'b0011100100011111; out_imag=16'b0001110011011101; end // in_theta = 0.148926 pi
 12'b000100110010: begin out_real=16'b0011100100010100; out_imag=16'b0001110011110011; end // in_theta = 0.149414 pi
 12'b000100110011: begin out_real=16'b0011100100001001; out_imag=16'b0001110100001010; end // in_theta = 0.149902 pi
 12'b000100110100: begin out_real=16'b0011100011111101; out_imag=16'b0001110100100000; end // in_theta = 0.150391 pi
 12'b000100110101: begin out_real=16'b0011100011110010; out_imag=16'b0001110100110110; end // in_theta = 0.150879 pi
 12'b000100110110: begin out_real=16'b0011100011100110; out_imag=16'b0001110101001101; end // in_theta = 0.151367 pi
 12'b000100110111: begin out_real=16'b0011100011011011; out_imag=16'b0001110101100011; end // in_theta = 0.151855 pi
 12'b000100111000: begin out_real=16'b0011100011001111; out_imag=16'b0001110101111001; end // in_theta = 0.152344 pi
 12'b000100111001: begin out_real=16'b0011100011000011; out_imag=16'b0001110110010000; end // in_theta = 0.152832 pi
 12'b000100111010: begin out_real=16'b0011100010111000; out_imag=16'b0001110110100110; end // in_theta = 0.153320 pi
 12'b000100111011: begin out_real=16'b0011100010101100; out_imag=16'b0001110110111100; end // in_theta = 0.153809 pi
 12'b000100111100: begin out_real=16'b0011100010100001; out_imag=16'b0001110111010011; end // in_theta = 0.154297 pi
 12'b000100111101: begin out_real=16'b0011100010010101; out_imag=16'b0001110111101001; end // in_theta = 0.154785 pi
 12'b000100111110: begin out_real=16'b0011100010001001; out_imag=16'b0001110111111111; end // in_theta = 0.155273 pi
 12'b000100111111: begin out_real=16'b0011100001111101; out_imag=16'b0001111000010101; end // in_theta = 0.155762 pi
 12'b000101000000: begin out_real=16'b0011100001110001; out_imag=16'b0001111000101011; end // in_theta = 0.156250 pi
 12'b000101000001: begin out_real=16'b0011100001100110; out_imag=16'b0001111001000010; end // in_theta = 0.156738 pi
 12'b000101000010: begin out_real=16'b0011100001011010; out_imag=16'b0001111001011000; end // in_theta = 0.157227 pi
 12'b000101000011: begin out_real=16'b0011100001001110; out_imag=16'b0001111001101110; end // in_theta = 0.157715 pi
 12'b000101000100: begin out_real=16'b0011100001000010; out_imag=16'b0001111010000100; end // in_theta = 0.158203 pi
 12'b000101000101: begin out_real=16'b0011100000110110; out_imag=16'b0001111010011010; end // in_theta = 0.158691 pi
 12'b000101000110: begin out_real=16'b0011100000101010; out_imag=16'b0001111010110000; end // in_theta = 0.159180 pi
 12'b000101000111: begin out_real=16'b0011100000011110; out_imag=16'b0001111011000110; end // in_theta = 0.159668 pi
 12'b000101001000: begin out_real=16'b0011100000010010; out_imag=16'b0001111011011100; end // in_theta = 0.160156 pi
 12'b000101001001: begin out_real=16'b0011100000000101; out_imag=16'b0001111011110010; end // in_theta = 0.160645 pi
 12'b000101001010: begin out_real=16'b0011011111111001; out_imag=16'b0001111100001000; end // in_theta = 0.161133 pi
 12'b000101001011: begin out_real=16'b0011011111101101; out_imag=16'b0001111100011110; end // in_theta = 0.161621 pi
 12'b000101001100: begin out_real=16'b0011011111100001; out_imag=16'b0001111100110100; end // in_theta = 0.162109 pi
 12'b000101001101: begin out_real=16'b0011011111010101; out_imag=16'b0001111101001010; end // in_theta = 0.162598 pi
 12'b000101001110: begin out_real=16'b0011011111001000; out_imag=16'b0001111101100000; end // in_theta = 0.163086 pi
 12'b000101001111: begin out_real=16'b0011011110111100; out_imag=16'b0001111101110110; end // in_theta = 0.163574 pi
 12'b000101010000: begin out_real=16'b0011011110110000; out_imag=16'b0001111110001100; end // in_theta = 0.164063 pi
 12'b000101010001: begin out_real=16'b0011011110100011; out_imag=16'b0001111110100010; end // in_theta = 0.164551 pi
 12'b000101010010: begin out_real=16'b0011011110010111; out_imag=16'b0001111110110111; end // in_theta = 0.165039 pi
 12'b000101010011: begin out_real=16'b0011011110001010; out_imag=16'b0001111111001101; end // in_theta = 0.165527 pi
 12'b000101010100: begin out_real=16'b0011011101111110; out_imag=16'b0001111111100011; end // in_theta = 0.166016 pi
 12'b000101010101: begin out_real=16'b0011011101110001; out_imag=16'b0001111111111001; end // in_theta = 0.166504 pi
 12'b000101010110: begin out_real=16'b0011011101100101; out_imag=16'b0010000000001111; end // in_theta = 0.166992 pi
 12'b000101010111: begin out_real=16'b0011011101011000; out_imag=16'b0010000000100100; end // in_theta = 0.167480 pi
 12'b000101011000: begin out_real=16'b0011011101001011; out_imag=16'b0010000000111010; end // in_theta = 0.167969 pi
 12'b000101011001: begin out_real=16'b0011011100111111; out_imag=16'b0010000001010000; end // in_theta = 0.168457 pi
 12'b000101011010: begin out_real=16'b0011011100110010; out_imag=16'b0010000001100101; end // in_theta = 0.168945 pi
 12'b000101011011: begin out_real=16'b0011011100100101; out_imag=16'b0010000001111011; end // in_theta = 0.169434 pi
 12'b000101011100: begin out_real=16'b0011011100011000; out_imag=16'b0010000010010001; end // in_theta = 0.169922 pi
 12'b000101011101: begin out_real=16'b0011011100001100; out_imag=16'b0010000010100110; end // in_theta = 0.170410 pi
 12'b000101011110: begin out_real=16'b0011011011111111; out_imag=16'b0010000010111100; end // in_theta = 0.170898 pi
 12'b000101011111: begin out_real=16'b0011011011110010; out_imag=16'b0010000011010001; end // in_theta = 0.171387 pi
 12'b000101100000: begin out_real=16'b0011011011100101; out_imag=16'b0010000011100111; end // in_theta = 0.171875 pi
 12'b000101100001: begin out_real=16'b0011011011011000; out_imag=16'b0010000011111101; end // in_theta = 0.172363 pi
 12'b000101100010: begin out_real=16'b0011011011001011; out_imag=16'b0010000100010010; end // in_theta = 0.172852 pi
 12'b000101100011: begin out_real=16'b0011011010111110; out_imag=16'b0010000100101000; end // in_theta = 0.173340 pi
 12'b000101100100: begin out_real=16'b0011011010110001; out_imag=16'b0010000100111101; end // in_theta = 0.173828 pi
 12'b000101100101: begin out_real=16'b0011011010100100; out_imag=16'b0010000101010011; end // in_theta = 0.174316 pi
 12'b000101100110: begin out_real=16'b0011011010010111; out_imag=16'b0010000101101000; end // in_theta = 0.174805 pi
 12'b000101100111: begin out_real=16'b0011011010001010; out_imag=16'b0010000101111101; end // in_theta = 0.175293 pi
 12'b000101101000: begin out_real=16'b0011011001111101; out_imag=16'b0010000110010011; end // in_theta = 0.175781 pi
 12'b000101101001: begin out_real=16'b0011011001101111; out_imag=16'b0010000110101000; end // in_theta = 0.176270 pi
 12'b000101101010: begin out_real=16'b0011011001100010; out_imag=16'b0010000110111110; end // in_theta = 0.176758 pi
 12'b000101101011: begin out_real=16'b0011011001010101; out_imag=16'b0010000111010011; end // in_theta = 0.177246 pi
 12'b000101101100: begin out_real=16'b0011011001001000; out_imag=16'b0010000111101000; end // in_theta = 0.177734 pi
 12'b000101101101: begin out_real=16'b0011011000111010; out_imag=16'b0010000111111110; end // in_theta = 0.178223 pi
 12'b000101101110: begin out_real=16'b0011011000101101; out_imag=16'b0010001000010011; end // in_theta = 0.178711 pi
 12'b000101101111: begin out_real=16'b0011011000100000; out_imag=16'b0010001000101000; end // in_theta = 0.179199 pi
 12'b000101110000: begin out_real=16'b0011011000010010; out_imag=16'b0010001000111101; end // in_theta = 0.179688 pi
 12'b000101110001: begin out_real=16'b0011011000000101; out_imag=16'b0010001001010011; end // in_theta = 0.180176 pi
 12'b000101110010: begin out_real=16'b0011010111110111; out_imag=16'b0010001001101000; end // in_theta = 0.180664 pi
 12'b000101110011: begin out_real=16'b0011010111101010; out_imag=16'b0010001001111101; end // in_theta = 0.181152 pi
 12'b000101110100: begin out_real=16'b0011010111011100; out_imag=16'b0010001010010010; end // in_theta = 0.181641 pi
 12'b000101110101: begin out_real=16'b0011010111001110; out_imag=16'b0010001010100111; end // in_theta = 0.182129 pi
 12'b000101110110: begin out_real=16'b0011010111000001; out_imag=16'b0010001010111100; end // in_theta = 0.182617 pi
 12'b000101110111: begin out_real=16'b0011010110110011; out_imag=16'b0010001011010010; end // in_theta = 0.183105 pi
 12'b000101111000: begin out_real=16'b0011010110100101; out_imag=16'b0010001011100111; end // in_theta = 0.183594 pi
 12'b000101111001: begin out_real=16'b0011010110011000; out_imag=16'b0010001011111100; end // in_theta = 0.184082 pi
 12'b000101111010: begin out_real=16'b0011010110001010; out_imag=16'b0010001100010001; end // in_theta = 0.184570 pi
 12'b000101111011: begin out_real=16'b0011010101111100; out_imag=16'b0010001100100110; end // in_theta = 0.185059 pi
 12'b000101111100: begin out_real=16'b0011010101101110; out_imag=16'b0010001100111011; end // in_theta = 0.185547 pi
 12'b000101111101: begin out_real=16'b0011010101100001; out_imag=16'b0010001101010000; end // in_theta = 0.186035 pi
 12'b000101111110: begin out_real=16'b0011010101010011; out_imag=16'b0010001101100101; end // in_theta = 0.186523 pi
 12'b000101111111: begin out_real=16'b0011010101000101; out_imag=16'b0010001101111010; end // in_theta = 0.187012 pi
 12'b000110000000: begin out_real=16'b0011010100110111; out_imag=16'b0010001110001110; end // in_theta = 0.187500 pi
 12'b000110000001: begin out_real=16'b0011010100101001; out_imag=16'b0010001110100011; end // in_theta = 0.187988 pi
 12'b000110000010: begin out_real=16'b0011010100011011; out_imag=16'b0010001110111000; end // in_theta = 0.188477 pi
 12'b000110000011: begin out_real=16'b0011010100001101; out_imag=16'b0010001111001101; end // in_theta = 0.188965 pi
 12'b000110000100: begin out_real=16'b0011010011111111; out_imag=16'b0010001111100010; end // in_theta = 0.189453 pi
 12'b000110000101: begin out_real=16'b0011010011110001; out_imag=16'b0010001111110111; end // in_theta = 0.189941 pi
 12'b000110000110: begin out_real=16'b0011010011100010; out_imag=16'b0010010000001011; end // in_theta = 0.190430 pi
 12'b000110000111: begin out_real=16'b0011010011010100; out_imag=16'b0010010000100000; end // in_theta = 0.190918 pi
 12'b000110001000: begin out_real=16'b0011010011000110; out_imag=16'b0010010000110101; end // in_theta = 0.191406 pi
 12'b000110001001: begin out_real=16'b0011010010111000; out_imag=16'b0010010001001010; end // in_theta = 0.191895 pi
 12'b000110001010: begin out_real=16'b0011010010101010; out_imag=16'b0010010001011110; end // in_theta = 0.192383 pi
 12'b000110001011: begin out_real=16'b0011010010011011; out_imag=16'b0010010001110011; end // in_theta = 0.192871 pi
 12'b000110001100: begin out_real=16'b0011010010001101; out_imag=16'b0010010010001000; end // in_theta = 0.193359 pi
 12'b000110001101: begin out_real=16'b0011010001111111; out_imag=16'b0010010010011100; end // in_theta = 0.193848 pi
 12'b000110001110: begin out_real=16'b0011010001110000; out_imag=16'b0010010010110001; end // in_theta = 0.194336 pi
 12'b000110001111: begin out_real=16'b0011010001100010; out_imag=16'b0010010011000101; end // in_theta = 0.194824 pi
 12'b000110010000: begin out_real=16'b0011010001010011; out_imag=16'b0010010011011010; end // in_theta = 0.195313 pi
 12'b000110010001: begin out_real=16'b0011010001000101; out_imag=16'b0010010011101111; end // in_theta = 0.195801 pi
 12'b000110010010: begin out_real=16'b0011010000110110; out_imag=16'b0010010100000011; end // in_theta = 0.196289 pi
 12'b000110010011: begin out_real=16'b0011010000101000; out_imag=16'b0010010100011000; end // in_theta = 0.196777 pi
 12'b000110010100: begin out_real=16'b0011010000011001; out_imag=16'b0010010100101100; end // in_theta = 0.197266 pi
 12'b000110010101: begin out_real=16'b0011010000001011; out_imag=16'b0010010101000001; end // in_theta = 0.197754 pi
 12'b000110010110: begin out_real=16'b0011001111111100; out_imag=16'b0010010101010101; end // in_theta = 0.198242 pi
 12'b000110010111: begin out_real=16'b0011001111101101; out_imag=16'b0010010101101001; end // in_theta = 0.198730 pi
 12'b000110011000: begin out_real=16'b0011001111011111; out_imag=16'b0010010101111110; end // in_theta = 0.199219 pi
 12'b000110011001: begin out_real=16'b0011001111010000; out_imag=16'b0010010110010010; end // in_theta = 0.199707 pi
 12'b000110011010: begin out_real=16'b0011001111000001; out_imag=16'b0010010110100110; end // in_theta = 0.200195 pi
 12'b000110011011: begin out_real=16'b0011001110110010; out_imag=16'b0010010110111011; end // in_theta = 0.200684 pi
 12'b000110011100: begin out_real=16'b0011001110100011; out_imag=16'b0010010111001111; end // in_theta = 0.201172 pi
 12'b000110011101: begin out_real=16'b0011001110010101; out_imag=16'b0010010111100011; end // in_theta = 0.201660 pi
 12'b000110011110: begin out_real=16'b0011001110000110; out_imag=16'b0010010111111000; end // in_theta = 0.202148 pi
 12'b000110011111: begin out_real=16'b0011001101110111; out_imag=16'b0010011000001100; end // in_theta = 0.202637 pi
 12'b000110100000: begin out_real=16'b0011001101101000; out_imag=16'b0010011000100000; end // in_theta = 0.203125 pi
 12'b000110100001: begin out_real=16'b0011001101011001; out_imag=16'b0010011000110100; end // in_theta = 0.203613 pi
 12'b000110100010: begin out_real=16'b0011001101001010; out_imag=16'b0010011001001000; end // in_theta = 0.204102 pi
 12'b000110100011: begin out_real=16'b0011001100111011; out_imag=16'b0010011001011100; end // in_theta = 0.204590 pi
 12'b000110100100: begin out_real=16'b0011001100101100; out_imag=16'b0010011001110001; end // in_theta = 0.205078 pi
 12'b000110100101: begin out_real=16'b0011001100011101; out_imag=16'b0010011010000101; end // in_theta = 0.205566 pi
 12'b000110100110: begin out_real=16'b0011001100001101; out_imag=16'b0010011010011001; end // in_theta = 0.206055 pi
 12'b000110100111: begin out_real=16'b0011001011111110; out_imag=16'b0010011010101101; end // in_theta = 0.206543 pi
 12'b000110101000: begin out_real=16'b0011001011101111; out_imag=16'b0010011011000001; end // in_theta = 0.207031 pi
 12'b000110101001: begin out_real=16'b0011001011100000; out_imag=16'b0010011011010101; end // in_theta = 0.207520 pi
 12'b000110101010: begin out_real=16'b0011001011010000; out_imag=16'b0010011011101001; end // in_theta = 0.208008 pi
 12'b000110101011: begin out_real=16'b0011001011000001; out_imag=16'b0010011011111101; end // in_theta = 0.208496 pi
 12'b000110101100: begin out_real=16'b0011001010110010; out_imag=16'b0010011100010001; end // in_theta = 0.208984 pi
 12'b000110101101: begin out_real=16'b0011001010100011; out_imag=16'b0010011100100100; end // in_theta = 0.209473 pi
 12'b000110101110: begin out_real=16'b0011001010010011; out_imag=16'b0010011100111000; end // in_theta = 0.209961 pi
 12'b000110101111: begin out_real=16'b0011001010000100; out_imag=16'b0010011101001100; end // in_theta = 0.210449 pi
 12'b000110110000: begin out_real=16'b0011001001110100; out_imag=16'b0010011101100000; end // in_theta = 0.210938 pi
 12'b000110110001: begin out_real=16'b0011001001100101; out_imag=16'b0010011101110100; end // in_theta = 0.211426 pi
 12'b000110110010: begin out_real=16'b0011001001010101; out_imag=16'b0010011110001000; end // in_theta = 0.211914 pi
 12'b000110110011: begin out_real=16'b0011001001000110; out_imag=16'b0010011110011011; end // in_theta = 0.212402 pi
 12'b000110110100: begin out_real=16'b0011001000110110; out_imag=16'b0010011110101111; end // in_theta = 0.212891 pi
 12'b000110110101: begin out_real=16'b0011001000100111; out_imag=16'b0010011111000011; end // in_theta = 0.213379 pi
 12'b000110110110: begin out_real=16'b0011001000010111; out_imag=16'b0010011111010110; end // in_theta = 0.213867 pi
 12'b000110110111: begin out_real=16'b0011001000000111; out_imag=16'b0010011111101010; end // in_theta = 0.214355 pi
 12'b000110111000: begin out_real=16'b0011000111111000; out_imag=16'b0010011111111110; end // in_theta = 0.214844 pi
 12'b000110111001: begin out_real=16'b0011000111101000; out_imag=16'b0010100000010001; end // in_theta = 0.215332 pi
 12'b000110111010: begin out_real=16'b0011000111011000; out_imag=16'b0010100000100101; end // in_theta = 0.215820 pi
 12'b000110111011: begin out_real=16'b0011000111001000; out_imag=16'b0010100000111000; end // in_theta = 0.216309 pi
 12'b000110111100: begin out_real=16'b0011000110111001; out_imag=16'b0010100001001100; end // in_theta = 0.216797 pi
 12'b000110111101: begin out_real=16'b0011000110101001; out_imag=16'b0010100001100000; end // in_theta = 0.217285 pi
 12'b000110111110: begin out_real=16'b0011000110011001; out_imag=16'b0010100001110011; end // in_theta = 0.217773 pi
 12'b000110111111: begin out_real=16'b0011000110001001; out_imag=16'b0010100010000110; end // in_theta = 0.218262 pi
 12'b000111000000: begin out_real=16'b0011000101111001; out_imag=16'b0010100010011010; end // in_theta = 0.218750 pi
 12'b000111000001: begin out_real=16'b0011000101101001; out_imag=16'b0010100010101101; end // in_theta = 0.219238 pi
 12'b000111000010: begin out_real=16'b0011000101011001; out_imag=16'b0010100011000001; end // in_theta = 0.219727 pi
 12'b000111000011: begin out_real=16'b0011000101001001; out_imag=16'b0010100011010100; end // in_theta = 0.220215 pi
 12'b000111000100: begin out_real=16'b0011000100111001; out_imag=16'b0010100011100111; end // in_theta = 0.220703 pi
 12'b000111000101: begin out_real=16'b0011000100101001; out_imag=16'b0010100011111011; end // in_theta = 0.221191 pi
 12'b000111000110: begin out_real=16'b0011000100011001; out_imag=16'b0010100100001110; end // in_theta = 0.221680 pi
 12'b000111000111: begin out_real=16'b0011000100001001; out_imag=16'b0010100100100001; end // in_theta = 0.222168 pi
 12'b000111001000: begin out_real=16'b0011000011111001; out_imag=16'b0010100100110101; end // in_theta = 0.222656 pi
 12'b000111001001: begin out_real=16'b0011000011101000; out_imag=16'b0010100101001000; end // in_theta = 0.223145 pi
 12'b000111001010: begin out_real=16'b0011000011011000; out_imag=16'b0010100101011011; end // in_theta = 0.223633 pi
 12'b000111001011: begin out_real=16'b0011000011001000; out_imag=16'b0010100101101110; end // in_theta = 0.224121 pi
 12'b000111001100: begin out_real=16'b0011000010111000; out_imag=16'b0010100110000001; end // in_theta = 0.224609 pi
 12'b000111001101: begin out_real=16'b0011000010100111; out_imag=16'b0010100110010100; end // in_theta = 0.225098 pi
 12'b000111001110: begin out_real=16'b0011000010010111; out_imag=16'b0010100110100111; end // in_theta = 0.225586 pi
 12'b000111001111: begin out_real=16'b0011000010000111; out_imag=16'b0010100110111011; end // in_theta = 0.226074 pi
 12'b000111010000: begin out_real=16'b0011000001110110; out_imag=16'b0010100111001110; end // in_theta = 0.226563 pi
 12'b000111010001: begin out_real=16'b0011000001100110; out_imag=16'b0010100111100001; end // in_theta = 0.227051 pi
 12'b000111010010: begin out_real=16'b0011000001010101; out_imag=16'b0010100111110100; end // in_theta = 0.227539 pi
 12'b000111010011: begin out_real=16'b0011000001000101; out_imag=16'b0010101000000111; end // in_theta = 0.228027 pi
 12'b000111010100: begin out_real=16'b0011000000110100; out_imag=16'b0010101000011010; end // in_theta = 0.228516 pi
 12'b000111010101: begin out_real=16'b0011000000100100; out_imag=16'b0010101000101100; end // in_theta = 0.229004 pi
 12'b000111010110: begin out_real=16'b0011000000010011; out_imag=16'b0010101000111111; end // in_theta = 0.229492 pi
 12'b000111010111: begin out_real=16'b0011000000000010; out_imag=16'b0010101001010010; end // in_theta = 0.229980 pi
 12'b000111011000: begin out_real=16'b0010111111110010; out_imag=16'b0010101001100101; end // in_theta = 0.230469 pi
 12'b000111011001: begin out_real=16'b0010111111100001; out_imag=16'b0010101001111000; end // in_theta = 0.230957 pi
 12'b000111011010: begin out_real=16'b0010111111010000; out_imag=16'b0010101010001011; end // in_theta = 0.231445 pi
 12'b000111011011: begin out_real=16'b0010111111000000; out_imag=16'b0010101010011101; end // in_theta = 0.231934 pi
 12'b000111011100: begin out_real=16'b0010111110101111; out_imag=16'b0010101010110000; end // in_theta = 0.232422 pi
 12'b000111011101: begin out_real=16'b0010111110011110; out_imag=16'b0010101011000011; end // in_theta = 0.232910 pi
 12'b000111011110: begin out_real=16'b0010111110001101; out_imag=16'b0010101011010110; end // in_theta = 0.233398 pi
 12'b000111011111: begin out_real=16'b0010111101111101; out_imag=16'b0010101011101000; end // in_theta = 0.233887 pi
 12'b000111100000: begin out_real=16'b0010111101101100; out_imag=16'b0010101011111011; end // in_theta = 0.234375 pi
 12'b000111100001: begin out_real=16'b0010111101011011; out_imag=16'b0010101100001101; end // in_theta = 0.234863 pi
 12'b000111100010: begin out_real=16'b0010111101001010; out_imag=16'b0010101100100000; end // in_theta = 0.235352 pi
 12'b000111100011: begin out_real=16'b0010111100111001; out_imag=16'b0010101100110011; end // in_theta = 0.235840 pi
 12'b000111100100: begin out_real=16'b0010111100101000; out_imag=16'b0010101101000101; end // in_theta = 0.236328 pi
 12'b000111100101: begin out_real=16'b0010111100010111; out_imag=16'b0010101101011000; end // in_theta = 0.236816 pi
 12'b000111100110: begin out_real=16'b0010111100000110; out_imag=16'b0010101101101010; end // in_theta = 0.237305 pi
 12'b000111100111: begin out_real=16'b0010111011110101; out_imag=16'b0010101101111101; end // in_theta = 0.237793 pi
 12'b000111101000: begin out_real=16'b0010111011100100; out_imag=16'b0010101110001111; end // in_theta = 0.238281 pi
 12'b000111101001: begin out_real=16'b0010111011010011; out_imag=16'b0010101110100001; end // in_theta = 0.238770 pi
 12'b000111101010: begin out_real=16'b0010111011000010; out_imag=16'b0010101110110100; end // in_theta = 0.239258 pi
 12'b000111101011: begin out_real=16'b0010111010110000; out_imag=16'b0010101111000110; end // in_theta = 0.239746 pi
 12'b000111101100: begin out_real=16'b0010111010011111; out_imag=16'b0010101111011000; end // in_theta = 0.240234 pi
 12'b000111101101: begin out_real=16'b0010111010001110; out_imag=16'b0010101111101011; end // in_theta = 0.240723 pi
 12'b000111101110: begin out_real=16'b0010111001111101; out_imag=16'b0010101111111101; end // in_theta = 0.241211 pi
 12'b000111101111: begin out_real=16'b0010111001101011; out_imag=16'b0010110000001111; end // in_theta = 0.241699 pi
 12'b000111110000: begin out_real=16'b0010111001011010; out_imag=16'b0010110000100001; end // in_theta = 0.242188 pi
 12'b000111110001: begin out_real=16'b0010111001001001; out_imag=16'b0010110000110100; end // in_theta = 0.242676 pi
 12'b000111110010: begin out_real=16'b0010111000110111; out_imag=16'b0010110001000110; end // in_theta = 0.243164 pi
 12'b000111110011: begin out_real=16'b0010111000100110; out_imag=16'b0010110001011000; end // in_theta = 0.243652 pi
 12'b000111110100: begin out_real=16'b0010111000010101; out_imag=16'b0010110001101010; end // in_theta = 0.244141 pi
 12'b000111110101: begin out_real=16'b0010111000000011; out_imag=16'b0010110001111100; end // in_theta = 0.244629 pi
 12'b000111110110: begin out_real=16'b0010110111110010; out_imag=16'b0010110010001110; end // in_theta = 0.245117 pi
 12'b000111110111: begin out_real=16'b0010110111100000; out_imag=16'b0010110010100000; end // in_theta = 0.245605 pi
 12'b000111111000: begin out_real=16'b0010110111001111; out_imag=16'b0010110010110010; end // in_theta = 0.246094 pi
 12'b000111111001: begin out_real=16'b0010110110111101; out_imag=16'b0010110011000100; end // in_theta = 0.246582 pi
 12'b000111111010: begin out_real=16'b0010110110101011; out_imag=16'b0010110011010110; end // in_theta = 0.247070 pi
 12'b000111111011: begin out_real=16'b0010110110011010; out_imag=16'b0010110011101000; end // in_theta = 0.247559 pi
 12'b000111111100: begin out_real=16'b0010110110001000; out_imag=16'b0010110011111010; end // in_theta = 0.248047 pi
 12'b000111111101: begin out_real=16'b0010110101110110; out_imag=16'b0010110100001100; end // in_theta = 0.248535 pi
 12'b000111111110: begin out_real=16'b0010110101100101; out_imag=16'b0010110100011110; end // in_theta = 0.249023 pi
 12'b000111111111: begin out_real=16'b0010110101010011; out_imag=16'b0010110100101111; end // in_theta = 0.249512 pi
 12'b001000000000: begin out_real=16'b0010110101000001; out_imag=16'b0010110101000001; end // in_theta = 0.250000 pi
 12'b001000000001: begin out_real=16'b0010110100101111; out_imag=16'b0010110101010011; end // in_theta = 0.250488 pi
 12'b001000000010: begin out_real=16'b0010110100011110; out_imag=16'b0010110101100101; end // in_theta = 0.250977 pi
 12'b001000000011: begin out_real=16'b0010110100001100; out_imag=16'b0010110101110110; end // in_theta = 0.251465 pi
 12'b001000000100: begin out_real=16'b0010110011111010; out_imag=16'b0010110110001000; end // in_theta = 0.251953 pi
 12'b001000000101: begin out_real=16'b0010110011101000; out_imag=16'b0010110110011010; end // in_theta = 0.252441 pi
 12'b001000000110: begin out_real=16'b0010110011010110; out_imag=16'b0010110110101011; end // in_theta = 0.252930 pi
 12'b001000000111: begin out_real=16'b0010110011000100; out_imag=16'b0010110110111101; end // in_theta = 0.253418 pi
 12'b001000001000: begin out_real=16'b0010110010110010; out_imag=16'b0010110111001111; end // in_theta = 0.253906 pi
 12'b001000001001: begin out_real=16'b0010110010100000; out_imag=16'b0010110111100000; end // in_theta = 0.254395 pi
 12'b001000001010: begin out_real=16'b0010110010001110; out_imag=16'b0010110111110010; end // in_theta = 0.254883 pi
 12'b001000001011: begin out_real=16'b0010110001111100; out_imag=16'b0010111000000011; end // in_theta = 0.255371 pi
 12'b001000001100: begin out_real=16'b0010110001101010; out_imag=16'b0010111000010101; end // in_theta = 0.255859 pi
 12'b001000001101: begin out_real=16'b0010110001011000; out_imag=16'b0010111000100110; end // in_theta = 0.256348 pi
 12'b001000001110: begin out_real=16'b0010110001000110; out_imag=16'b0010111000110111; end // in_theta = 0.256836 pi
 12'b001000001111: begin out_real=16'b0010110000110100; out_imag=16'b0010111001001001; end // in_theta = 0.257324 pi
 12'b001000010000: begin out_real=16'b0010110000100001; out_imag=16'b0010111001011010; end // in_theta = 0.257813 pi
 12'b001000010001: begin out_real=16'b0010110000001111; out_imag=16'b0010111001101011; end // in_theta = 0.258301 pi
 12'b001000010010: begin out_real=16'b0010101111111101; out_imag=16'b0010111001111101; end // in_theta = 0.258789 pi
 12'b001000010011: begin out_real=16'b0010101111101011; out_imag=16'b0010111010001110; end // in_theta = 0.259277 pi
 12'b001000010100: begin out_real=16'b0010101111011000; out_imag=16'b0010111010011111; end // in_theta = 0.259766 pi
 12'b001000010101: begin out_real=16'b0010101111000110; out_imag=16'b0010111010110000; end // in_theta = 0.260254 pi
 12'b001000010110: begin out_real=16'b0010101110110100; out_imag=16'b0010111011000010; end // in_theta = 0.260742 pi
 12'b001000010111: begin out_real=16'b0010101110100001; out_imag=16'b0010111011010011; end // in_theta = 0.261230 pi
 12'b001000011000: begin out_real=16'b0010101110001111; out_imag=16'b0010111011100100; end // in_theta = 0.261719 pi
 12'b001000011001: begin out_real=16'b0010101101111101; out_imag=16'b0010111011110101; end // in_theta = 0.262207 pi
 12'b001000011010: begin out_real=16'b0010101101101010; out_imag=16'b0010111100000110; end // in_theta = 0.262695 pi
 12'b001000011011: begin out_real=16'b0010101101011000; out_imag=16'b0010111100010111; end // in_theta = 0.263184 pi
 12'b001000011100: begin out_real=16'b0010101101000101; out_imag=16'b0010111100101000; end // in_theta = 0.263672 pi
 12'b001000011101: begin out_real=16'b0010101100110011; out_imag=16'b0010111100111001; end // in_theta = 0.264160 pi
 12'b001000011110: begin out_real=16'b0010101100100000; out_imag=16'b0010111101001010; end // in_theta = 0.264648 pi
 12'b001000011111: begin out_real=16'b0010101100001101; out_imag=16'b0010111101011011; end // in_theta = 0.265137 pi
 12'b001000100000: begin out_real=16'b0010101011111011; out_imag=16'b0010111101101100; end // in_theta = 0.265625 pi
 12'b001000100001: begin out_real=16'b0010101011101000; out_imag=16'b0010111101111101; end // in_theta = 0.266113 pi
 12'b001000100010: begin out_real=16'b0010101011010110; out_imag=16'b0010111110001101; end // in_theta = 0.266602 pi
 12'b001000100011: begin out_real=16'b0010101011000011; out_imag=16'b0010111110011110; end // in_theta = 0.267090 pi
 12'b001000100100: begin out_real=16'b0010101010110000; out_imag=16'b0010111110101111; end // in_theta = 0.267578 pi
 12'b001000100101: begin out_real=16'b0010101010011101; out_imag=16'b0010111111000000; end // in_theta = 0.268066 pi
 12'b001000100110: begin out_real=16'b0010101010001011; out_imag=16'b0010111111010000; end // in_theta = 0.268555 pi
 12'b001000100111: begin out_real=16'b0010101001111000; out_imag=16'b0010111111100001; end // in_theta = 0.269043 pi
 12'b001000101000: begin out_real=16'b0010101001100101; out_imag=16'b0010111111110010; end // in_theta = 0.269531 pi
 12'b001000101001: begin out_real=16'b0010101001010010; out_imag=16'b0011000000000010; end // in_theta = 0.270020 pi
 12'b001000101010: begin out_real=16'b0010101000111111; out_imag=16'b0011000000010011; end // in_theta = 0.270508 pi
 12'b001000101011: begin out_real=16'b0010101000101100; out_imag=16'b0011000000100100; end // in_theta = 0.270996 pi
 12'b001000101100: begin out_real=16'b0010101000011010; out_imag=16'b0011000000110100; end // in_theta = 0.271484 pi
 12'b001000101101: begin out_real=16'b0010101000000111; out_imag=16'b0011000001000101; end // in_theta = 0.271973 pi
 12'b001000101110: begin out_real=16'b0010100111110100; out_imag=16'b0011000001010101; end // in_theta = 0.272461 pi
 12'b001000101111: begin out_real=16'b0010100111100001; out_imag=16'b0011000001100110; end // in_theta = 0.272949 pi
 12'b001000110000: begin out_real=16'b0010100111001110; out_imag=16'b0011000001110110; end // in_theta = 0.273438 pi
 12'b001000110001: begin out_real=16'b0010100110111011; out_imag=16'b0011000010000111; end // in_theta = 0.273926 pi
 12'b001000110010: begin out_real=16'b0010100110100111; out_imag=16'b0011000010010111; end // in_theta = 0.274414 pi
 12'b001000110011: begin out_real=16'b0010100110010100; out_imag=16'b0011000010100111; end // in_theta = 0.274902 pi
 12'b001000110100: begin out_real=16'b0010100110000001; out_imag=16'b0011000010111000; end // in_theta = 0.275391 pi
 12'b001000110101: begin out_real=16'b0010100101101110; out_imag=16'b0011000011001000; end // in_theta = 0.275879 pi
 12'b001000110110: begin out_real=16'b0010100101011011; out_imag=16'b0011000011011000; end // in_theta = 0.276367 pi
 12'b001000110111: begin out_real=16'b0010100101001000; out_imag=16'b0011000011101000; end // in_theta = 0.276855 pi
 12'b001000111000: begin out_real=16'b0010100100110101; out_imag=16'b0011000011111001; end // in_theta = 0.277344 pi
 12'b001000111001: begin out_real=16'b0010100100100001; out_imag=16'b0011000100001001; end // in_theta = 0.277832 pi
 12'b001000111010: begin out_real=16'b0010100100001110; out_imag=16'b0011000100011001; end // in_theta = 0.278320 pi
 12'b001000111011: begin out_real=16'b0010100011111011; out_imag=16'b0011000100101001; end // in_theta = 0.278809 pi
 12'b001000111100: begin out_real=16'b0010100011100111; out_imag=16'b0011000100111001; end // in_theta = 0.279297 pi
 12'b001000111101: begin out_real=16'b0010100011010100; out_imag=16'b0011000101001001; end // in_theta = 0.279785 pi
 12'b001000111110: begin out_real=16'b0010100011000001; out_imag=16'b0011000101011001; end // in_theta = 0.280273 pi
 12'b001000111111: begin out_real=16'b0010100010101101; out_imag=16'b0011000101101001; end // in_theta = 0.280762 pi
 12'b001001000000: begin out_real=16'b0010100010011010; out_imag=16'b0011000101111001; end // in_theta = 0.281250 pi
 12'b001001000001: begin out_real=16'b0010100010000110; out_imag=16'b0011000110001001; end // in_theta = 0.281738 pi
 12'b001001000010: begin out_real=16'b0010100001110011; out_imag=16'b0011000110011001; end // in_theta = 0.282227 pi
 12'b001001000011: begin out_real=16'b0010100001100000; out_imag=16'b0011000110101001; end // in_theta = 0.282715 pi
 12'b001001000100: begin out_real=16'b0010100001001100; out_imag=16'b0011000110111001; end // in_theta = 0.283203 pi
 12'b001001000101: begin out_real=16'b0010100000111000; out_imag=16'b0011000111001000; end // in_theta = 0.283691 pi
 12'b001001000110: begin out_real=16'b0010100000100101; out_imag=16'b0011000111011000; end // in_theta = 0.284180 pi
 12'b001001000111: begin out_real=16'b0010100000010001; out_imag=16'b0011000111101000; end // in_theta = 0.284668 pi
 12'b001001001000: begin out_real=16'b0010011111111110; out_imag=16'b0011000111111000; end // in_theta = 0.285156 pi
 12'b001001001001: begin out_real=16'b0010011111101010; out_imag=16'b0011001000000111; end // in_theta = 0.285645 pi
 12'b001001001010: begin out_real=16'b0010011111010110; out_imag=16'b0011001000010111; end // in_theta = 0.286133 pi
 12'b001001001011: begin out_real=16'b0010011111000011; out_imag=16'b0011001000100111; end // in_theta = 0.286621 pi
 12'b001001001100: begin out_real=16'b0010011110101111; out_imag=16'b0011001000110110; end // in_theta = 0.287109 pi
 12'b001001001101: begin out_real=16'b0010011110011011; out_imag=16'b0011001001000110; end // in_theta = 0.287598 pi
 12'b001001001110: begin out_real=16'b0010011110001000; out_imag=16'b0011001001010101; end // in_theta = 0.288086 pi
 12'b001001001111: begin out_real=16'b0010011101110100; out_imag=16'b0011001001100101; end // in_theta = 0.288574 pi
 12'b001001010000: begin out_real=16'b0010011101100000; out_imag=16'b0011001001110100; end // in_theta = 0.289063 pi
 12'b001001010001: begin out_real=16'b0010011101001100; out_imag=16'b0011001010000100; end // in_theta = 0.289551 pi
 12'b001001010010: begin out_real=16'b0010011100111000; out_imag=16'b0011001010010011; end // in_theta = 0.290039 pi
 12'b001001010011: begin out_real=16'b0010011100100100; out_imag=16'b0011001010100011; end // in_theta = 0.290527 pi
 12'b001001010100: begin out_real=16'b0010011100010001; out_imag=16'b0011001010110010; end // in_theta = 0.291016 pi
 12'b001001010101: begin out_real=16'b0010011011111101; out_imag=16'b0011001011000001; end // in_theta = 0.291504 pi
 12'b001001010110: begin out_real=16'b0010011011101001; out_imag=16'b0011001011010000; end // in_theta = 0.291992 pi
 12'b001001010111: begin out_real=16'b0010011011010101; out_imag=16'b0011001011100000; end // in_theta = 0.292480 pi
 12'b001001011000: begin out_real=16'b0010011011000001; out_imag=16'b0011001011101111; end // in_theta = 0.292969 pi
 12'b001001011001: begin out_real=16'b0010011010101101; out_imag=16'b0011001011111110; end // in_theta = 0.293457 pi
 12'b001001011010: begin out_real=16'b0010011010011001; out_imag=16'b0011001100001101; end // in_theta = 0.293945 pi
 12'b001001011011: begin out_real=16'b0010011010000101; out_imag=16'b0011001100011101; end // in_theta = 0.294434 pi
 12'b001001011100: begin out_real=16'b0010011001110001; out_imag=16'b0011001100101100; end // in_theta = 0.294922 pi
 12'b001001011101: begin out_real=16'b0010011001011100; out_imag=16'b0011001100111011; end // in_theta = 0.295410 pi
 12'b001001011110: begin out_real=16'b0010011001001000; out_imag=16'b0011001101001010; end // in_theta = 0.295898 pi
 12'b001001011111: begin out_real=16'b0010011000110100; out_imag=16'b0011001101011001; end // in_theta = 0.296387 pi
 12'b001001100000: begin out_real=16'b0010011000100000; out_imag=16'b0011001101101000; end // in_theta = 0.296875 pi
 12'b001001100001: begin out_real=16'b0010011000001100; out_imag=16'b0011001101110111; end // in_theta = 0.297363 pi
 12'b001001100010: begin out_real=16'b0010010111111000; out_imag=16'b0011001110000110; end // in_theta = 0.297852 pi
 12'b001001100011: begin out_real=16'b0010010111100011; out_imag=16'b0011001110010101; end // in_theta = 0.298340 pi
 12'b001001100100: begin out_real=16'b0010010111001111; out_imag=16'b0011001110100011; end // in_theta = 0.298828 pi
 12'b001001100101: begin out_real=16'b0010010110111011; out_imag=16'b0011001110110010; end // in_theta = 0.299316 pi
 12'b001001100110: begin out_real=16'b0010010110100110; out_imag=16'b0011001111000001; end // in_theta = 0.299805 pi
 12'b001001100111: begin out_real=16'b0010010110010010; out_imag=16'b0011001111010000; end // in_theta = 0.300293 pi
 12'b001001101000: begin out_real=16'b0010010101111110; out_imag=16'b0011001111011111; end // in_theta = 0.300781 pi
 12'b001001101001: begin out_real=16'b0010010101101001; out_imag=16'b0011001111101101; end // in_theta = 0.301270 pi
 12'b001001101010: begin out_real=16'b0010010101010101; out_imag=16'b0011001111111100; end // in_theta = 0.301758 pi
 12'b001001101011: begin out_real=16'b0010010101000001; out_imag=16'b0011010000001011; end // in_theta = 0.302246 pi
 12'b001001101100: begin out_real=16'b0010010100101100; out_imag=16'b0011010000011001; end // in_theta = 0.302734 pi
 12'b001001101101: begin out_real=16'b0010010100011000; out_imag=16'b0011010000101000; end // in_theta = 0.303223 pi
 12'b001001101110: begin out_real=16'b0010010100000011; out_imag=16'b0011010000110110; end // in_theta = 0.303711 pi
 12'b001001101111: begin out_real=16'b0010010011101111; out_imag=16'b0011010001000101; end // in_theta = 0.304199 pi
 12'b001001110000: begin out_real=16'b0010010011011010; out_imag=16'b0011010001010011; end // in_theta = 0.304688 pi
 12'b001001110001: begin out_real=16'b0010010011000101; out_imag=16'b0011010001100010; end // in_theta = 0.305176 pi
 12'b001001110010: begin out_real=16'b0010010010110001; out_imag=16'b0011010001110000; end // in_theta = 0.305664 pi
 12'b001001110011: begin out_real=16'b0010010010011100; out_imag=16'b0011010001111111; end // in_theta = 0.306152 pi
 12'b001001110100: begin out_real=16'b0010010010001000; out_imag=16'b0011010010001101; end // in_theta = 0.306641 pi
 12'b001001110101: begin out_real=16'b0010010001110011; out_imag=16'b0011010010011011; end // in_theta = 0.307129 pi
 12'b001001110110: begin out_real=16'b0010010001011110; out_imag=16'b0011010010101010; end // in_theta = 0.307617 pi
 12'b001001110111: begin out_real=16'b0010010001001010; out_imag=16'b0011010010111000; end // in_theta = 0.308105 pi
 12'b001001111000: begin out_real=16'b0010010000110101; out_imag=16'b0011010011000110; end // in_theta = 0.308594 pi
 12'b001001111001: begin out_real=16'b0010010000100000; out_imag=16'b0011010011010100; end // in_theta = 0.309082 pi
 12'b001001111010: begin out_real=16'b0010010000001011; out_imag=16'b0011010011100010; end // in_theta = 0.309570 pi
 12'b001001111011: begin out_real=16'b0010001111110111; out_imag=16'b0011010011110001; end // in_theta = 0.310059 pi
 12'b001001111100: begin out_real=16'b0010001111100010; out_imag=16'b0011010011111111; end // in_theta = 0.310547 pi
 12'b001001111101: begin out_real=16'b0010001111001101; out_imag=16'b0011010100001101; end // in_theta = 0.311035 pi
 12'b001001111110: begin out_real=16'b0010001110111000; out_imag=16'b0011010100011011; end // in_theta = 0.311523 pi
 12'b001001111111: begin out_real=16'b0010001110100011; out_imag=16'b0011010100101001; end // in_theta = 0.312012 pi
 12'b001010000000: begin out_real=16'b0010001110001110; out_imag=16'b0011010100110111; end // in_theta = 0.312500 pi
 12'b001010000001: begin out_real=16'b0010001101111010; out_imag=16'b0011010101000101; end // in_theta = 0.312988 pi
 12'b001010000010: begin out_real=16'b0010001101100101; out_imag=16'b0011010101010011; end // in_theta = 0.313477 pi
 12'b001010000011: begin out_real=16'b0010001101010000; out_imag=16'b0011010101100001; end // in_theta = 0.313965 pi
 12'b001010000100: begin out_real=16'b0010001100111011; out_imag=16'b0011010101101110; end // in_theta = 0.314453 pi
 12'b001010000101: begin out_real=16'b0010001100100110; out_imag=16'b0011010101111100; end // in_theta = 0.314941 pi
 12'b001010000110: begin out_real=16'b0010001100010001; out_imag=16'b0011010110001010; end // in_theta = 0.315430 pi
 12'b001010000111: begin out_real=16'b0010001011111100; out_imag=16'b0011010110011000; end // in_theta = 0.315918 pi
 12'b001010001000: begin out_real=16'b0010001011100111; out_imag=16'b0011010110100101; end // in_theta = 0.316406 pi
 12'b001010001001: begin out_real=16'b0010001011010010; out_imag=16'b0011010110110011; end // in_theta = 0.316895 pi
 12'b001010001010: begin out_real=16'b0010001010111100; out_imag=16'b0011010111000001; end // in_theta = 0.317383 pi
 12'b001010001011: begin out_real=16'b0010001010100111; out_imag=16'b0011010111001110; end // in_theta = 0.317871 pi
 12'b001010001100: begin out_real=16'b0010001010010010; out_imag=16'b0011010111011100; end // in_theta = 0.318359 pi
 12'b001010001101: begin out_real=16'b0010001001111101; out_imag=16'b0011010111101010; end // in_theta = 0.318848 pi
 12'b001010001110: begin out_real=16'b0010001001101000; out_imag=16'b0011010111110111; end // in_theta = 0.319336 pi
 12'b001010001111: begin out_real=16'b0010001001010011; out_imag=16'b0011011000000101; end // in_theta = 0.319824 pi
 12'b001010010000: begin out_real=16'b0010001000111101; out_imag=16'b0011011000010010; end // in_theta = 0.320313 pi
 12'b001010010001: begin out_real=16'b0010001000101000; out_imag=16'b0011011000100000; end // in_theta = 0.320801 pi
 12'b001010010010: begin out_real=16'b0010001000010011; out_imag=16'b0011011000101101; end // in_theta = 0.321289 pi
 12'b001010010011: begin out_real=16'b0010000111111110; out_imag=16'b0011011000111010; end // in_theta = 0.321777 pi
 12'b001010010100: begin out_real=16'b0010000111101000; out_imag=16'b0011011001001000; end // in_theta = 0.322266 pi
 12'b001010010101: begin out_real=16'b0010000111010011; out_imag=16'b0011011001010101; end // in_theta = 0.322754 pi
 12'b001010010110: begin out_real=16'b0010000110111110; out_imag=16'b0011011001100010; end // in_theta = 0.323242 pi
 12'b001010010111: begin out_real=16'b0010000110101000; out_imag=16'b0011011001101111; end // in_theta = 0.323730 pi
 12'b001010011000: begin out_real=16'b0010000110010011; out_imag=16'b0011011001111101; end // in_theta = 0.324219 pi
 12'b001010011001: begin out_real=16'b0010000101111101; out_imag=16'b0011011010001010; end // in_theta = 0.324707 pi
 12'b001010011010: begin out_real=16'b0010000101101000; out_imag=16'b0011011010010111; end // in_theta = 0.325195 pi
 12'b001010011011: begin out_real=16'b0010000101010011; out_imag=16'b0011011010100100; end // in_theta = 0.325684 pi
 12'b001010011100: begin out_real=16'b0010000100111101; out_imag=16'b0011011010110001; end // in_theta = 0.326172 pi
 12'b001010011101: begin out_real=16'b0010000100101000; out_imag=16'b0011011010111110; end // in_theta = 0.326660 pi
 12'b001010011110: begin out_real=16'b0010000100010010; out_imag=16'b0011011011001011; end // in_theta = 0.327148 pi
 12'b001010011111: begin out_real=16'b0010000011111101; out_imag=16'b0011011011011000; end // in_theta = 0.327637 pi
 12'b001010100000: begin out_real=16'b0010000011100111; out_imag=16'b0011011011100101; end // in_theta = 0.328125 pi
 12'b001010100001: begin out_real=16'b0010000011010001; out_imag=16'b0011011011110010; end // in_theta = 0.328613 pi
 12'b001010100010: begin out_real=16'b0010000010111100; out_imag=16'b0011011011111111; end // in_theta = 0.329102 pi
 12'b001010100011: begin out_real=16'b0010000010100110; out_imag=16'b0011011100001100; end // in_theta = 0.329590 pi
 12'b001010100100: begin out_real=16'b0010000010010001; out_imag=16'b0011011100011000; end // in_theta = 0.330078 pi
 12'b001010100101: begin out_real=16'b0010000001111011; out_imag=16'b0011011100100101; end // in_theta = 0.330566 pi
 12'b001010100110: begin out_real=16'b0010000001100101; out_imag=16'b0011011100110010; end // in_theta = 0.331055 pi
 12'b001010100111: begin out_real=16'b0010000001010000; out_imag=16'b0011011100111111; end // in_theta = 0.331543 pi
 12'b001010101000: begin out_real=16'b0010000000111010; out_imag=16'b0011011101001011; end // in_theta = 0.332031 pi
 12'b001010101001: begin out_real=16'b0010000000100100; out_imag=16'b0011011101011000; end // in_theta = 0.332520 pi
 12'b001010101010: begin out_real=16'b0010000000001111; out_imag=16'b0011011101100101; end // in_theta = 0.333008 pi
 12'b001010101011: begin out_real=16'b0001111111111001; out_imag=16'b0011011101110001; end // in_theta = 0.333496 pi
 12'b001010101100: begin out_real=16'b0001111111100011; out_imag=16'b0011011101111110; end // in_theta = 0.333984 pi
 12'b001010101101: begin out_real=16'b0001111111001101; out_imag=16'b0011011110001010; end // in_theta = 0.334473 pi
 12'b001010101110: begin out_real=16'b0001111110110111; out_imag=16'b0011011110010111; end // in_theta = 0.334961 pi
 12'b001010101111: begin out_real=16'b0001111110100010; out_imag=16'b0011011110100011; end // in_theta = 0.335449 pi
 12'b001010110000: begin out_real=16'b0001111110001100; out_imag=16'b0011011110110000; end // in_theta = 0.335938 pi
 12'b001010110001: begin out_real=16'b0001111101110110; out_imag=16'b0011011110111100; end // in_theta = 0.336426 pi
 12'b001010110010: begin out_real=16'b0001111101100000; out_imag=16'b0011011111001000; end // in_theta = 0.336914 pi
 12'b001010110011: begin out_real=16'b0001111101001010; out_imag=16'b0011011111010101; end // in_theta = 0.337402 pi
 12'b001010110100: begin out_real=16'b0001111100110100; out_imag=16'b0011011111100001; end // in_theta = 0.337891 pi
 12'b001010110101: begin out_real=16'b0001111100011110; out_imag=16'b0011011111101101; end // in_theta = 0.338379 pi
 12'b001010110110: begin out_real=16'b0001111100001000; out_imag=16'b0011011111111001; end // in_theta = 0.338867 pi
 12'b001010110111: begin out_real=16'b0001111011110010; out_imag=16'b0011100000000101; end // in_theta = 0.339355 pi
 12'b001010111000: begin out_real=16'b0001111011011100; out_imag=16'b0011100000010010; end // in_theta = 0.339844 pi
 12'b001010111001: begin out_real=16'b0001111011000110; out_imag=16'b0011100000011110; end // in_theta = 0.340332 pi
 12'b001010111010: begin out_real=16'b0001111010110000; out_imag=16'b0011100000101010; end // in_theta = 0.340820 pi
 12'b001010111011: begin out_real=16'b0001111010011010; out_imag=16'b0011100000110110; end // in_theta = 0.341309 pi
 12'b001010111100: begin out_real=16'b0001111010000100; out_imag=16'b0011100001000010; end // in_theta = 0.341797 pi
 12'b001010111101: begin out_real=16'b0001111001101110; out_imag=16'b0011100001001110; end // in_theta = 0.342285 pi
 12'b001010111110: begin out_real=16'b0001111001011000; out_imag=16'b0011100001011010; end // in_theta = 0.342773 pi
 12'b001010111111: begin out_real=16'b0001111001000010; out_imag=16'b0011100001100110; end // in_theta = 0.343262 pi
 12'b001011000000: begin out_real=16'b0001111000101011; out_imag=16'b0011100001110001; end // in_theta = 0.343750 pi
 12'b001011000001: begin out_real=16'b0001111000010101; out_imag=16'b0011100001111101; end // in_theta = 0.344238 pi
 12'b001011000010: begin out_real=16'b0001110111111111; out_imag=16'b0011100010001001; end // in_theta = 0.344727 pi
 12'b001011000011: begin out_real=16'b0001110111101001; out_imag=16'b0011100010010101; end // in_theta = 0.345215 pi
 12'b001011000100: begin out_real=16'b0001110111010011; out_imag=16'b0011100010100001; end // in_theta = 0.345703 pi
 12'b001011000101: begin out_real=16'b0001110110111100; out_imag=16'b0011100010101100; end // in_theta = 0.346191 pi
 12'b001011000110: begin out_real=16'b0001110110100110; out_imag=16'b0011100010111000; end // in_theta = 0.346680 pi
 12'b001011000111: begin out_real=16'b0001110110010000; out_imag=16'b0011100011000011; end // in_theta = 0.347168 pi
 12'b001011001000: begin out_real=16'b0001110101111001; out_imag=16'b0011100011001111; end // in_theta = 0.347656 pi
 12'b001011001001: begin out_real=16'b0001110101100011; out_imag=16'b0011100011011011; end // in_theta = 0.348145 pi
 12'b001011001010: begin out_real=16'b0001110101001101; out_imag=16'b0011100011100110; end // in_theta = 0.348633 pi
 12'b001011001011: begin out_real=16'b0001110100110110; out_imag=16'b0011100011110010; end // in_theta = 0.349121 pi
 12'b001011001100: begin out_real=16'b0001110100100000; out_imag=16'b0011100011111101; end // in_theta = 0.349609 pi
 12'b001011001101: begin out_real=16'b0001110100001010; out_imag=16'b0011100100001001; end // in_theta = 0.350098 pi
 12'b001011001110: begin out_real=16'b0001110011110011; out_imag=16'b0011100100010100; end // in_theta = 0.350586 pi
 12'b001011001111: begin out_real=16'b0001110011011101; out_imag=16'b0011100100011111; end // in_theta = 0.351074 pi
 12'b001011010000: begin out_real=16'b0001110011000110; out_imag=16'b0011100100101011; end // in_theta = 0.351563 pi
 12'b001011010001: begin out_real=16'b0001110010110000; out_imag=16'b0011100100110110; end // in_theta = 0.352051 pi
 12'b001011010010: begin out_real=16'b0001110010011001; out_imag=16'b0011100101000001; end // in_theta = 0.352539 pi
 12'b001011010011: begin out_real=16'b0001110010000011; out_imag=16'b0011100101001100; end // in_theta = 0.353027 pi
 12'b001011010100: begin out_real=16'b0001110001101100; out_imag=16'b0011100101011000; end // in_theta = 0.353516 pi
 12'b001011010101: begin out_real=16'b0001110001010110; out_imag=16'b0011100101100011; end // in_theta = 0.354004 pi
 12'b001011010110: begin out_real=16'b0001110000111111; out_imag=16'b0011100101101110; end // in_theta = 0.354492 pi
 12'b001011010111: begin out_real=16'b0001110000101001; out_imag=16'b0011100101111001; end // in_theta = 0.354980 pi
 12'b001011011000: begin out_real=16'b0001110000010010; out_imag=16'b0011100110000100; end // in_theta = 0.355469 pi
 12'b001011011001: begin out_real=16'b0001101111111100; out_imag=16'b0011100110001111; end // in_theta = 0.355957 pi
 12'b001011011010: begin out_real=16'b0001101111100101; out_imag=16'b0011100110011010; end // in_theta = 0.356445 pi
 12'b001011011011: begin out_real=16'b0001101111001110; out_imag=16'b0011100110100101; end // in_theta = 0.356934 pi
 12'b001011011100: begin out_real=16'b0001101110111000; out_imag=16'b0011100110110000; end // in_theta = 0.357422 pi
 12'b001011011101: begin out_real=16'b0001101110100001; out_imag=16'b0011100110111011; end // in_theta = 0.357910 pi
 12'b001011011110: begin out_real=16'b0001101110001010; out_imag=16'b0011100111000101; end // in_theta = 0.358398 pi
 12'b001011011111: begin out_real=16'b0001101101110100; out_imag=16'b0011100111010000; end // in_theta = 0.358887 pi
 12'b001011100000: begin out_real=16'b0001101101011101; out_imag=16'b0011100111011011; end // in_theta = 0.359375 pi
 12'b001011100001: begin out_real=16'b0001101101000110; out_imag=16'b0011100111100110; end // in_theta = 0.359863 pi
 12'b001011100010: begin out_real=16'b0001101100110000; out_imag=16'b0011100111110000; end // in_theta = 0.360352 pi
 12'b001011100011: begin out_real=16'b0001101100011001; out_imag=16'b0011100111111011; end // in_theta = 0.360840 pi
 12'b001011100100: begin out_real=16'b0001101100000010; out_imag=16'b0011101000000110; end // in_theta = 0.361328 pi
 12'b001011100101: begin out_real=16'b0001101011101011; out_imag=16'b0011101000010000; end // in_theta = 0.361816 pi
 12'b001011100110: begin out_real=16'b0001101011010100; out_imag=16'b0011101000011011; end // in_theta = 0.362305 pi
 12'b001011100111: begin out_real=16'b0001101010111110; out_imag=16'b0011101000100101; end // in_theta = 0.362793 pi
 12'b001011101000: begin out_real=16'b0001101010100111; out_imag=16'b0011101000110000; end // in_theta = 0.363281 pi
 12'b001011101001: begin out_real=16'b0001101010010000; out_imag=16'b0011101000111010; end // in_theta = 0.363770 pi
 12'b001011101010: begin out_real=16'b0001101001111001; out_imag=16'b0011101001000101; end // in_theta = 0.364258 pi
 12'b001011101011: begin out_real=16'b0001101001100010; out_imag=16'b0011101001001111; end // in_theta = 0.364746 pi
 12'b001011101100: begin out_real=16'b0001101001001011; out_imag=16'b0011101001011001; end // in_theta = 0.365234 pi
 12'b001011101101: begin out_real=16'b0001101000110100; out_imag=16'b0011101001100100; end // in_theta = 0.365723 pi
 12'b001011101110: begin out_real=16'b0001101000011101; out_imag=16'b0011101001101110; end // in_theta = 0.366211 pi
 12'b001011101111: begin out_real=16'b0001101000000110; out_imag=16'b0011101001111000; end // in_theta = 0.366699 pi
 12'b001011110000: begin out_real=16'b0001100111101111; out_imag=16'b0011101010000010; end // in_theta = 0.367188 pi
 12'b001011110001: begin out_real=16'b0001100111011000; out_imag=16'b0011101010001101; end // in_theta = 0.367676 pi
 12'b001011110010: begin out_real=16'b0001100111000001; out_imag=16'b0011101010010111; end // in_theta = 0.368164 pi
 12'b001011110011: begin out_real=16'b0001100110101010; out_imag=16'b0011101010100001; end // in_theta = 0.368652 pi
 12'b001011110100: begin out_real=16'b0001100110010011; out_imag=16'b0011101010101011; end // in_theta = 0.369141 pi
 12'b001011110101: begin out_real=16'b0001100101111100; out_imag=16'b0011101010110101; end // in_theta = 0.369629 pi
 12'b001011110110: begin out_real=16'b0001100101100101; out_imag=16'b0011101010111111; end // in_theta = 0.370117 pi
 12'b001011110111: begin out_real=16'b0001100101001110; out_imag=16'b0011101011001001; end // in_theta = 0.370605 pi
 12'b001011111000: begin out_real=16'b0001100100110111; out_imag=16'b0011101011010011; end // in_theta = 0.371094 pi
 12'b001011111001: begin out_real=16'b0001100100100000; out_imag=16'b0011101011011101; end // in_theta = 0.371582 pi
 12'b001011111010: begin out_real=16'b0001100100001001; out_imag=16'b0011101011100110; end // in_theta = 0.372070 pi
 12'b001011111011: begin out_real=16'b0001100011110010; out_imag=16'b0011101011110000; end // in_theta = 0.372559 pi
 12'b001011111100: begin out_real=16'b0001100011011011; out_imag=16'b0011101011111010; end // in_theta = 0.373047 pi
 12'b001011111101: begin out_real=16'b0001100011000011; out_imag=16'b0011101100000100; end // in_theta = 0.373535 pi
 12'b001011111110: begin out_real=16'b0001100010101100; out_imag=16'b0011101100001110; end // in_theta = 0.374023 pi
 12'b001011111111: begin out_real=16'b0001100010010101; out_imag=16'b0011101100010111; end // in_theta = 0.374512 pi
 12'b001100000000: begin out_real=16'b0001100001111110; out_imag=16'b0011101100100001; end // in_theta = 0.375000 pi
 12'b001100000001: begin out_real=16'b0001100001100111; out_imag=16'b0011101100101010; end // in_theta = 0.375488 pi
 12'b001100000010: begin out_real=16'b0001100001001111; out_imag=16'b0011101100110100; end // in_theta = 0.375977 pi
 12'b001100000011: begin out_real=16'b0001100000111000; out_imag=16'b0011101100111110; end // in_theta = 0.376465 pi
 12'b001100000100: begin out_real=16'b0001100000100001; out_imag=16'b0011101101000111; end // in_theta = 0.376953 pi
 12'b001100000101: begin out_real=16'b0001100000001010; out_imag=16'b0011101101010000; end // in_theta = 0.377441 pi
 12'b001100000110: begin out_real=16'b0001011111110010; out_imag=16'b0011101101011010; end // in_theta = 0.377930 pi
 12'b001100000111: begin out_real=16'b0001011111011011; out_imag=16'b0011101101100011; end // in_theta = 0.378418 pi
 12'b001100001000: begin out_real=16'b0001011111000100; out_imag=16'b0011101101101101; end // in_theta = 0.378906 pi
 12'b001100001001: begin out_real=16'b0001011110101100; out_imag=16'b0011101101110110; end // in_theta = 0.379395 pi
 12'b001100001010: begin out_real=16'b0001011110010101; out_imag=16'b0011101101111111; end // in_theta = 0.379883 pi
 12'b001100001011: begin out_real=16'b0001011101111110; out_imag=16'b0011101110001000; end // in_theta = 0.380371 pi
 12'b001100001100: begin out_real=16'b0001011101100110; out_imag=16'b0011101110010010; end // in_theta = 0.380859 pi
 12'b001100001101: begin out_real=16'b0001011101001111; out_imag=16'b0011101110011011; end // in_theta = 0.381348 pi
 12'b001100001110: begin out_real=16'b0001011100110111; out_imag=16'b0011101110100100; end // in_theta = 0.381836 pi
 12'b001100001111: begin out_real=16'b0001011100100000; out_imag=16'b0011101110101101; end // in_theta = 0.382324 pi
 12'b001100010000: begin out_real=16'b0001011100001001; out_imag=16'b0011101110110110; end // in_theta = 0.382813 pi
 12'b001100010001: begin out_real=16'b0001011011110001; out_imag=16'b0011101110111111; end // in_theta = 0.383301 pi
 12'b001100010010: begin out_real=16'b0001011011011010; out_imag=16'b0011101111001000; end // in_theta = 0.383789 pi
 12'b001100010011: begin out_real=16'b0001011011000010; out_imag=16'b0011101111010001; end // in_theta = 0.384277 pi
 12'b001100010100: begin out_real=16'b0001011010101011; out_imag=16'b0011101111011010; end // in_theta = 0.384766 pi
 12'b001100010101: begin out_real=16'b0001011010010011; out_imag=16'b0011101111100011; end // in_theta = 0.385254 pi
 12'b001100010110: begin out_real=16'b0001011001111100; out_imag=16'b0011101111101100; end // in_theta = 0.385742 pi
 12'b001100010111: begin out_real=16'b0001011001100100; out_imag=16'b0011101111110101; end // in_theta = 0.386230 pi
 12'b001100011000: begin out_real=16'b0001011001001100; out_imag=16'b0011101111111101; end // in_theta = 0.386719 pi
 12'b001100011001: begin out_real=16'b0001011000110101; out_imag=16'b0011110000000110; end // in_theta = 0.387207 pi
 12'b001100011010: begin out_real=16'b0001011000011101; out_imag=16'b0011110000001111; end // in_theta = 0.387695 pi
 12'b001100011011: begin out_real=16'b0001011000000110; out_imag=16'b0011110000010111; end // in_theta = 0.388184 pi
 12'b001100011100: begin out_real=16'b0001010111101110; out_imag=16'b0011110000100000; end // in_theta = 0.388672 pi
 12'b001100011101: begin out_real=16'b0001010111010111; out_imag=16'b0011110000101001; end // in_theta = 0.389160 pi
 12'b001100011110: begin out_real=16'b0001010110111111; out_imag=16'b0011110000110001; end // in_theta = 0.389648 pi
 12'b001100011111: begin out_real=16'b0001010110100111; out_imag=16'b0011110000111010; end // in_theta = 0.390137 pi
 12'b001100100000: begin out_real=16'b0001010110010000; out_imag=16'b0011110001000010; end // in_theta = 0.390625 pi
 12'b001100100001: begin out_real=16'b0001010101111000; out_imag=16'b0011110001001011; end // in_theta = 0.391113 pi
 12'b001100100010: begin out_real=16'b0001010101100000; out_imag=16'b0011110001010011; end // in_theta = 0.391602 pi
 12'b001100100011: begin out_real=16'b0001010101001001; out_imag=16'b0011110001011011; end // in_theta = 0.392090 pi
 12'b001100100100: begin out_real=16'b0001010100110001; out_imag=16'b0011110001100100; end // in_theta = 0.392578 pi
 12'b001100100101: begin out_real=16'b0001010100011001; out_imag=16'b0011110001101100; end // in_theta = 0.393066 pi
 12'b001100100110: begin out_real=16'b0001010100000001; out_imag=16'b0011110001110100; end // in_theta = 0.393555 pi
 12'b001100100111: begin out_real=16'b0001010011101010; out_imag=16'b0011110001111101; end // in_theta = 0.394043 pi
 12'b001100101000: begin out_real=16'b0001010011010010; out_imag=16'b0011110010000101; end // in_theta = 0.394531 pi
 12'b001100101001: begin out_real=16'b0001010010111010; out_imag=16'b0011110010001101; end // in_theta = 0.395020 pi
 12'b001100101010: begin out_real=16'b0001010010100010; out_imag=16'b0011110010010101; end // in_theta = 0.395508 pi
 12'b001100101011: begin out_real=16'b0001010010001011; out_imag=16'b0011110010011101; end // in_theta = 0.395996 pi
 12'b001100101100: begin out_real=16'b0001010001110011; out_imag=16'b0011110010100101; end // in_theta = 0.396484 pi
 12'b001100101101: begin out_real=16'b0001010001011011; out_imag=16'b0011110010101101; end // in_theta = 0.396973 pi
 12'b001100101110: begin out_real=16'b0001010001000011; out_imag=16'b0011110010110101; end // in_theta = 0.397461 pi
 12'b001100101111: begin out_real=16'b0001010000101011; out_imag=16'b0011110010111101; end // in_theta = 0.397949 pi
 12'b001100110000: begin out_real=16'b0001010000010011; out_imag=16'b0011110011000101; end // in_theta = 0.398438 pi
 12'b001100110001: begin out_real=16'b0001001111111011; out_imag=16'b0011110011001101; end // in_theta = 0.398926 pi
 12'b001100110010: begin out_real=16'b0001001111100100; out_imag=16'b0011110011010101; end // in_theta = 0.399414 pi
 12'b001100110011: begin out_real=16'b0001001111001100; out_imag=16'b0011110011011101; end // in_theta = 0.399902 pi
 12'b001100110100: begin out_real=16'b0001001110110100; out_imag=16'b0011110011100100; end // in_theta = 0.400391 pi
 12'b001100110101: begin out_real=16'b0001001110011100; out_imag=16'b0011110011101100; end // in_theta = 0.400879 pi
 12'b001100110110: begin out_real=16'b0001001110000100; out_imag=16'b0011110011110100; end // in_theta = 0.401367 pi
 12'b001100110111: begin out_real=16'b0001001101101100; out_imag=16'b0011110011111011; end // in_theta = 0.401855 pi
 12'b001100111000: begin out_real=16'b0001001101010100; out_imag=16'b0011110100000011; end // in_theta = 0.402344 pi
 12'b001100111001: begin out_real=16'b0001001100111100; out_imag=16'b0011110100001011; end // in_theta = 0.402832 pi
 12'b001100111010: begin out_real=16'b0001001100100100; out_imag=16'b0011110100010010; end // in_theta = 0.403320 pi
 12'b001100111011: begin out_real=16'b0001001100001100; out_imag=16'b0011110100011010; end // in_theta = 0.403809 pi
 12'b001100111100: begin out_real=16'b0001001011110100; out_imag=16'b0011110100100001; end // in_theta = 0.404297 pi
 12'b001100111101: begin out_real=16'b0001001011011100; out_imag=16'b0011110100101000; end // in_theta = 0.404785 pi
 12'b001100111110: begin out_real=16'b0001001011000100; out_imag=16'b0011110100110000; end // in_theta = 0.405273 pi
 12'b001100111111: begin out_real=16'b0001001010101100; out_imag=16'b0011110100110111; end // in_theta = 0.405762 pi
 12'b001101000000: begin out_real=16'b0001001010010100; out_imag=16'b0011110100111111; end // in_theta = 0.406250 pi
 12'b001101000001: begin out_real=16'b0001001001111100; out_imag=16'b0011110101000110; end // in_theta = 0.406738 pi
 12'b001101000010: begin out_real=16'b0001001001100100; out_imag=16'b0011110101001101; end // in_theta = 0.407227 pi
 12'b001101000011: begin out_real=16'b0001001001001100; out_imag=16'b0011110101010100; end // in_theta = 0.407715 pi
 12'b001101000100: begin out_real=16'b0001001000110100; out_imag=16'b0011110101011011; end // in_theta = 0.408203 pi
 12'b001101000101: begin out_real=16'b0001001000011100; out_imag=16'b0011110101100011; end // in_theta = 0.408691 pi
 12'b001101000110: begin out_real=16'b0001001000000100; out_imag=16'b0011110101101010; end // in_theta = 0.409180 pi
 12'b001101000111: begin out_real=16'b0001000111101011; out_imag=16'b0011110101110001; end // in_theta = 0.409668 pi
 12'b001101001000: begin out_real=16'b0001000111010011; out_imag=16'b0011110101111000; end // in_theta = 0.410156 pi
 12'b001101001001: begin out_real=16'b0001000110111011; out_imag=16'b0011110101111111; end // in_theta = 0.410645 pi
 12'b001101001010: begin out_real=16'b0001000110100011; out_imag=16'b0011110110000110; end // in_theta = 0.411133 pi
 12'b001101001011: begin out_real=16'b0001000110001011; out_imag=16'b0011110110001101; end // in_theta = 0.411621 pi
 12'b001101001100: begin out_real=16'b0001000101110011; out_imag=16'b0011110110010011; end // in_theta = 0.412109 pi
 12'b001101001101: begin out_real=16'b0001000101011010; out_imag=16'b0011110110011010; end // in_theta = 0.412598 pi
 12'b001101001110: begin out_real=16'b0001000101000010; out_imag=16'b0011110110100001; end // in_theta = 0.413086 pi
 12'b001101001111: begin out_real=16'b0001000100101010; out_imag=16'b0011110110101000; end // in_theta = 0.413574 pi
 12'b001101010000: begin out_real=16'b0001000100010010; out_imag=16'b0011110110101111; end // in_theta = 0.414063 pi
 12'b001101010001: begin out_real=16'b0001000011111010; out_imag=16'b0011110110110101; end // in_theta = 0.414551 pi
 12'b001101010010: begin out_real=16'b0001000011100001; out_imag=16'b0011110110111100; end // in_theta = 0.415039 pi
 12'b001101010011: begin out_real=16'b0001000011001001; out_imag=16'b0011110111000010; end // in_theta = 0.415527 pi
 12'b001101010100: begin out_real=16'b0001000010110001; out_imag=16'b0011110111001001; end // in_theta = 0.416016 pi
 12'b001101010101: begin out_real=16'b0001000010011001; out_imag=16'b0011110111010000; end // in_theta = 0.416504 pi
 12'b001101010110: begin out_real=16'b0001000010000000; out_imag=16'b0011110111010110; end // in_theta = 0.416992 pi
 12'b001101010111: begin out_real=16'b0001000001101000; out_imag=16'b0011110111011101; end // in_theta = 0.417480 pi
 12'b001101011000: begin out_real=16'b0001000001010000; out_imag=16'b0011110111100011; end // in_theta = 0.417969 pi
 12'b001101011001: begin out_real=16'b0001000000110111; out_imag=16'b0011110111101001; end // in_theta = 0.418457 pi
 12'b001101011010: begin out_real=16'b0001000000011111; out_imag=16'b0011110111110000; end // in_theta = 0.418945 pi
 12'b001101011011: begin out_real=16'b0001000000000111; out_imag=16'b0011110111110110; end // in_theta = 0.419434 pi
 12'b001101011100: begin out_real=16'b0000111111101110; out_imag=16'b0011110111111100; end // in_theta = 0.419922 pi
 12'b001101011101: begin out_real=16'b0000111111010110; out_imag=16'b0011111000000011; end // in_theta = 0.420410 pi
 12'b001101011110: begin out_real=16'b0000111110111110; out_imag=16'b0011111000001001; end // in_theta = 0.420898 pi
 12'b001101011111: begin out_real=16'b0000111110100101; out_imag=16'b0011111000001111; end // in_theta = 0.421387 pi
 12'b001101100000: begin out_real=16'b0000111110001101; out_imag=16'b0011111000010101; end // in_theta = 0.421875 pi
 12'b001101100001: begin out_real=16'b0000111101110101; out_imag=16'b0011111000011011; end // in_theta = 0.422363 pi
 12'b001101100010: begin out_real=16'b0000111101011100; out_imag=16'b0011111000100001; end // in_theta = 0.422852 pi
 12'b001101100011: begin out_real=16'b0000111101000100; out_imag=16'b0011111000100111; end // in_theta = 0.423340 pi
 12'b001101100100: begin out_real=16'b0000111100101011; out_imag=16'b0011111000101101; end // in_theta = 0.423828 pi
 12'b001101100101: begin out_real=16'b0000111100010011; out_imag=16'b0011111000110011; end // in_theta = 0.424316 pi
 12'b001101100110: begin out_real=16'b0000111011111011; out_imag=16'b0011111000111001; end // in_theta = 0.424805 pi
 12'b001101100111: begin out_real=16'b0000111011100010; out_imag=16'b0011111000111111; end // in_theta = 0.425293 pi
 12'b001101101000: begin out_real=16'b0000111011001010; out_imag=16'b0011111001000101; end // in_theta = 0.425781 pi
 12'b001101101001: begin out_real=16'b0000111010110001; out_imag=16'b0011111001001010; end // in_theta = 0.426270 pi
 12'b001101101010: begin out_real=16'b0000111010011001; out_imag=16'b0011111001010000; end // in_theta = 0.426758 pi
 12'b001101101011: begin out_real=16'b0000111010000000; out_imag=16'b0011111001010110; end // in_theta = 0.427246 pi
 12'b001101101100: begin out_real=16'b0000111001101000; out_imag=16'b0011111001011100; end // in_theta = 0.427734 pi
 12'b001101101101: begin out_real=16'b0000111001001111; out_imag=16'b0011111001100001; end // in_theta = 0.428223 pi
 12'b001101101110: begin out_real=16'b0000111000110111; out_imag=16'b0011111001100111; end // in_theta = 0.428711 pi
 12'b001101101111: begin out_real=16'b0000111000011110; out_imag=16'b0011111001101100; end // in_theta = 0.429199 pi
 12'b001101110000: begin out_real=16'b0000111000000110; out_imag=16'b0011111001110010; end // in_theta = 0.429688 pi
 12'b001101110001: begin out_real=16'b0000110111101101; out_imag=16'b0011111001110111; end // in_theta = 0.430176 pi
 12'b001101110010: begin out_real=16'b0000110111010101; out_imag=16'b0011111001111101; end // in_theta = 0.430664 pi
 12'b001101110011: begin out_real=16'b0000110110111100; out_imag=16'b0011111010000010; end // in_theta = 0.431152 pi
 12'b001101110100: begin out_real=16'b0000110110100100; out_imag=16'b0011111010001000; end // in_theta = 0.431641 pi
 12'b001101110101: begin out_real=16'b0000110110001011; out_imag=16'b0011111010001101; end // in_theta = 0.432129 pi
 12'b001101110110: begin out_real=16'b0000110101110010; out_imag=16'b0011111010010010; end // in_theta = 0.432617 pi
 12'b001101110111: begin out_real=16'b0000110101011010; out_imag=16'b0011111010011000; end // in_theta = 0.433105 pi
 12'b001101111000: begin out_real=16'b0000110101000001; out_imag=16'b0011111010011101; end // in_theta = 0.433594 pi
 12'b001101111001: begin out_real=16'b0000110100101001; out_imag=16'b0011111010100010; end // in_theta = 0.434082 pi
 12'b001101111010: begin out_real=16'b0000110100010000; out_imag=16'b0011111010100111; end // in_theta = 0.434570 pi
 12'b001101111011: begin out_real=16'b0000110011111000; out_imag=16'b0011111010101100; end // in_theta = 0.435059 pi
 12'b001101111100: begin out_real=16'b0000110011011111; out_imag=16'b0011111010110001; end // in_theta = 0.435547 pi
 12'b001101111101: begin out_real=16'b0000110011000110; out_imag=16'b0011111010110110; end // in_theta = 0.436035 pi
 12'b001101111110: begin out_real=16'b0000110010101110; out_imag=16'b0011111010111011; end // in_theta = 0.436523 pi
 12'b001101111111: begin out_real=16'b0000110010010101; out_imag=16'b0011111011000000; end // in_theta = 0.437012 pi
 12'b001110000000: begin out_real=16'b0000110001111100; out_imag=16'b0011111011000101; end // in_theta = 0.437500 pi
 12'b001110000001: begin out_real=16'b0000110001100100; out_imag=16'b0011111011001010; end // in_theta = 0.437988 pi
 12'b001110000010: begin out_real=16'b0000110001001011; out_imag=16'b0011111011001111; end // in_theta = 0.438477 pi
 12'b001110000011: begin out_real=16'b0000110000110010; out_imag=16'b0011111011010100; end // in_theta = 0.438965 pi
 12'b001110000100: begin out_real=16'b0000110000011010; out_imag=16'b0011111011011000; end // in_theta = 0.439453 pi
 12'b001110000101: begin out_real=16'b0000110000000001; out_imag=16'b0011111011011101; end // in_theta = 0.439941 pi
 12'b001110000110: begin out_real=16'b0000101111101000; out_imag=16'b0011111011100010; end // in_theta = 0.440430 pi
 12'b001110000111: begin out_real=16'b0000101111010000; out_imag=16'b0011111011100111; end // in_theta = 0.440918 pi
 12'b001110001000: begin out_real=16'b0000101110110111; out_imag=16'b0011111011101011; end // in_theta = 0.441406 pi
 12'b001110001001: begin out_real=16'b0000101110011110; out_imag=16'b0011111011110000; end // in_theta = 0.441895 pi
 12'b001110001010: begin out_real=16'b0000101110000101; out_imag=16'b0011111011110100; end // in_theta = 0.442383 pi
 12'b001110001011: begin out_real=16'b0000101101101101; out_imag=16'b0011111011111001; end // in_theta = 0.442871 pi
 12'b001110001100: begin out_real=16'b0000101101010100; out_imag=16'b0011111011111101; end // in_theta = 0.443359 pi
 12'b001110001101: begin out_real=16'b0000101100111011; out_imag=16'b0011111100000010; end // in_theta = 0.443848 pi
 12'b001110001110: begin out_real=16'b0000101100100011; out_imag=16'b0011111100000110; end // in_theta = 0.444336 pi
 12'b001110001111: begin out_real=16'b0000101100001010; out_imag=16'b0011111100001010; end // in_theta = 0.444824 pi
 12'b001110010000: begin out_real=16'b0000101011110001; out_imag=16'b0011111100001111; end // in_theta = 0.445313 pi
 12'b001110010001: begin out_real=16'b0000101011011000; out_imag=16'b0011111100010011; end // in_theta = 0.445801 pi
 12'b001110010010: begin out_real=16'b0000101011000000; out_imag=16'b0011111100010111; end // in_theta = 0.446289 pi
 12'b001110010011: begin out_real=16'b0000101010100111; out_imag=16'b0011111100011100; end // in_theta = 0.446777 pi
 12'b001110010100: begin out_real=16'b0000101010001110; out_imag=16'b0011111100100000; end // in_theta = 0.447266 pi
 12'b001110010101: begin out_real=16'b0000101001110101; out_imag=16'b0011111100100100; end // in_theta = 0.447754 pi
 12'b001110010110: begin out_real=16'b0000101001011100; out_imag=16'b0011111100101000; end // in_theta = 0.448242 pi
 12'b001110010111: begin out_real=16'b0000101001000100; out_imag=16'b0011111100101100; end // in_theta = 0.448730 pi
 12'b001110011000: begin out_real=16'b0000101000101011; out_imag=16'b0011111100110000; end // in_theta = 0.449219 pi
 12'b001110011001: begin out_real=16'b0000101000010010; out_imag=16'b0011111100110100; end // in_theta = 0.449707 pi
 12'b001110011010: begin out_real=16'b0000100111111001; out_imag=16'b0011111100111000; end // in_theta = 0.450195 pi
 12'b001110011011: begin out_real=16'b0000100111100000; out_imag=16'b0011111100111100; end // in_theta = 0.450684 pi
 12'b001110011100: begin out_real=16'b0000100111000111; out_imag=16'b0011111101000000; end // in_theta = 0.451172 pi
 12'b001110011101: begin out_real=16'b0000100110101111; out_imag=16'b0011111101000011; end // in_theta = 0.451660 pi
 12'b001110011110: begin out_real=16'b0000100110010110; out_imag=16'b0011111101000111; end // in_theta = 0.452148 pi
 12'b001110011111: begin out_real=16'b0000100101111101; out_imag=16'b0011111101001011; end // in_theta = 0.452637 pi
 12'b001110100000: begin out_real=16'b0000100101100100; out_imag=16'b0011111101001111; end // in_theta = 0.453125 pi
 12'b001110100001: begin out_real=16'b0000100101001011; out_imag=16'b0011111101010010; end // in_theta = 0.453613 pi
 12'b001110100010: begin out_real=16'b0000100100110010; out_imag=16'b0011111101010110; end // in_theta = 0.454102 pi
 12'b001110100011: begin out_real=16'b0000100100011001; out_imag=16'b0011111101011010; end // in_theta = 0.454590 pi
 12'b001110100100: begin out_real=16'b0000100100000001; out_imag=16'b0011111101011101; end // in_theta = 0.455078 pi
 12'b001110100101: begin out_real=16'b0000100011101000; out_imag=16'b0011111101100001; end // in_theta = 0.455566 pi
 12'b001110100110: begin out_real=16'b0000100011001111; out_imag=16'b0011111101100100; end // in_theta = 0.456055 pi
 12'b001110100111: begin out_real=16'b0000100010110110; out_imag=16'b0011111101101000; end // in_theta = 0.456543 pi
 12'b001110101000: begin out_real=16'b0000100010011101; out_imag=16'b0011111101101011; end // in_theta = 0.457031 pi
 12'b001110101001: begin out_real=16'b0000100010000100; out_imag=16'b0011111101101110; end // in_theta = 0.457520 pi
 12'b001110101010: begin out_real=16'b0000100001101011; out_imag=16'b0011111101110010; end // in_theta = 0.458008 pi
 12'b001110101011: begin out_real=16'b0000100001010010; out_imag=16'b0011111101110101; end // in_theta = 0.458496 pi
 12'b001110101100: begin out_real=16'b0000100000111001; out_imag=16'b0011111101111000; end // in_theta = 0.458984 pi
 12'b001110101101: begin out_real=16'b0000100000100000; out_imag=16'b0011111101111011; end // in_theta = 0.459473 pi
 12'b001110101110: begin out_real=16'b0000100000000111; out_imag=16'b0011111101111111; end // in_theta = 0.459961 pi
 12'b001110101111: begin out_real=16'b0000011111101111; out_imag=16'b0011111110000010; end // in_theta = 0.460449 pi
 12'b001110110000: begin out_real=16'b0000011111010110; out_imag=16'b0011111110000101; end // in_theta = 0.460938 pi
 12'b001110110001: begin out_real=16'b0000011110111101; out_imag=16'b0011111110001000; end // in_theta = 0.461426 pi
 12'b001110110010: begin out_real=16'b0000011110100100; out_imag=16'b0011111110001011; end // in_theta = 0.461914 pi
 12'b001110110011: begin out_real=16'b0000011110001011; out_imag=16'b0011111110001110; end // in_theta = 0.462402 pi
 12'b001110110100: begin out_real=16'b0000011101110010; out_imag=16'b0011111110010001; end // in_theta = 0.462891 pi
 12'b001110110101: begin out_real=16'b0000011101011001; out_imag=16'b0011111110010100; end // in_theta = 0.463379 pi
 12'b001110110110: begin out_real=16'b0000011101000000; out_imag=16'b0011111110010111; end // in_theta = 0.463867 pi
 12'b001110110111: begin out_real=16'b0000011100100111; out_imag=16'b0011111110011001; end // in_theta = 0.464355 pi
 12'b001110111000: begin out_real=16'b0000011100001110; out_imag=16'b0011111110011100; end // in_theta = 0.464844 pi
 12'b001110111001: begin out_real=16'b0000011011110101; out_imag=16'b0011111110011111; end // in_theta = 0.465332 pi
 12'b001110111010: begin out_real=16'b0000011011011100; out_imag=16'b0011111110100010; end // in_theta = 0.465820 pi
 12'b001110111011: begin out_real=16'b0000011011000011; out_imag=16'b0011111110100100; end // in_theta = 0.466309 pi
 12'b001110111100: begin out_real=16'b0000011010101010; out_imag=16'b0011111110100111; end // in_theta = 0.466797 pi
 12'b001110111101: begin out_real=16'b0000011010010001; out_imag=16'b0011111110101010; end // in_theta = 0.467285 pi
 12'b001110111110: begin out_real=16'b0000011001111000; out_imag=16'b0011111110101100; end // in_theta = 0.467773 pi
 12'b001110111111: begin out_real=16'b0000011001011111; out_imag=16'b0011111110101111; end // in_theta = 0.468262 pi
 12'b001111000000: begin out_real=16'b0000011001000110; out_imag=16'b0011111110110001; end // in_theta = 0.468750 pi
 12'b001111000001: begin out_real=16'b0000011000101101; out_imag=16'b0011111110110100; end // in_theta = 0.469238 pi
 12'b001111000010: begin out_real=16'b0000011000010100; out_imag=16'b0011111110110110; end // in_theta = 0.469727 pi
 12'b001111000011: begin out_real=16'b0000010111111011; out_imag=16'b0011111110111000; end // in_theta = 0.470215 pi
 12'b001111000100: begin out_real=16'b0000010111100010; out_imag=16'b0011111110111011; end // in_theta = 0.470703 pi
 12'b001111000101: begin out_real=16'b0000010111001001; out_imag=16'b0011111110111101; end // in_theta = 0.471191 pi
 12'b001111000110: begin out_real=16'b0000010110110000; out_imag=16'b0011111110111111; end // in_theta = 0.471680 pi
 12'b001111000111: begin out_real=16'b0000010110010111; out_imag=16'b0011111111000001; end // in_theta = 0.472168 pi
 12'b001111001000: begin out_real=16'b0000010101111110; out_imag=16'b0011111111000100; end // in_theta = 0.472656 pi
 12'b001111001001: begin out_real=16'b0000010101100101; out_imag=16'b0011111111000110; end // in_theta = 0.473145 pi
 12'b001111001010: begin out_real=16'b0000010101001100; out_imag=16'b0011111111001000; end // in_theta = 0.473633 pi
 12'b001111001011: begin out_real=16'b0000010100110011; out_imag=16'b0011111111001010; end // in_theta = 0.474121 pi
 12'b001111001100: begin out_real=16'b0000010100011010; out_imag=16'b0011111111001100; end // in_theta = 0.474609 pi
 12'b001111001101: begin out_real=16'b0000010100000000; out_imag=16'b0011111111001110; end // in_theta = 0.475098 pi
 12'b001111001110: begin out_real=16'b0000010011100111; out_imag=16'b0011111111010000; end // in_theta = 0.475586 pi
 12'b001111001111: begin out_real=16'b0000010011001110; out_imag=16'b0011111111010010; end // in_theta = 0.476074 pi
 12'b001111010000: begin out_real=16'b0000010010110101; out_imag=16'b0011111111010100; end // in_theta = 0.476563 pi
 12'b001111010001: begin out_real=16'b0000010010011100; out_imag=16'b0011111111010101; end // in_theta = 0.477051 pi
 12'b001111010010: begin out_real=16'b0000010010000011; out_imag=16'b0011111111010111; end // in_theta = 0.477539 pi
 12'b001111010011: begin out_real=16'b0000010001101010; out_imag=16'b0011111111011001; end // in_theta = 0.478027 pi
 12'b001111010100: begin out_real=16'b0000010001010001; out_imag=16'b0011111111011011; end // in_theta = 0.478516 pi
 12'b001111010101: begin out_real=16'b0000010000111000; out_imag=16'b0011111111011100; end // in_theta = 0.479004 pi
 12'b001111010110: begin out_real=16'b0000010000011111; out_imag=16'b0011111111011110; end // in_theta = 0.479492 pi
 12'b001111010111: begin out_real=16'b0000010000000110; out_imag=16'b0011111111100000; end // in_theta = 0.479980 pi
 12'b001111011000: begin out_real=16'b0000001111101101; out_imag=16'b0011111111100001; end // in_theta = 0.480469 pi
 12'b001111011001: begin out_real=16'b0000001111010100; out_imag=16'b0011111111100011; end // in_theta = 0.480957 pi
 12'b001111011010: begin out_real=16'b0000001110111011; out_imag=16'b0011111111100100; end // in_theta = 0.481445 pi
 12'b001111011011: begin out_real=16'b0000001110100001; out_imag=16'b0011111111100110; end // in_theta = 0.481934 pi
 12'b001111011100: begin out_real=16'b0000001110001000; out_imag=16'b0011111111100111; end // in_theta = 0.482422 pi
 12'b001111011101: begin out_real=16'b0000001101101111; out_imag=16'b0011111111101000; end // in_theta = 0.482910 pi
 12'b001111011110: begin out_real=16'b0000001101010110; out_imag=16'b0011111111101010; end // in_theta = 0.483398 pi
 12'b001111011111: begin out_real=16'b0000001100111101; out_imag=16'b0011111111101011; end // in_theta = 0.483887 pi
 12'b001111100000: begin out_real=16'b0000001100100100; out_imag=16'b0011111111101100; end // in_theta = 0.484375 pi
 12'b001111100001: begin out_real=16'b0000001100001011; out_imag=16'b0011111111101101; end // in_theta = 0.484863 pi
 12'b001111100010: begin out_real=16'b0000001011110010; out_imag=16'b0011111111101111; end // in_theta = 0.485352 pi
 12'b001111100011: begin out_real=16'b0000001011011001; out_imag=16'b0011111111110000; end // in_theta = 0.485840 pi
 12'b001111100100: begin out_real=16'b0000001011000000; out_imag=16'b0011111111110001; end // in_theta = 0.486328 pi
 12'b001111100101: begin out_real=16'b0000001010100110; out_imag=16'b0011111111110010; end // in_theta = 0.486816 pi
 12'b001111100110: begin out_real=16'b0000001010001101; out_imag=16'b0011111111110011; end // in_theta = 0.487305 pi
 12'b001111100111: begin out_real=16'b0000001001110100; out_imag=16'b0011111111110100; end // in_theta = 0.487793 pi
 12'b001111101000: begin out_real=16'b0000001001011011; out_imag=16'b0011111111110101; end // in_theta = 0.488281 pi
 12'b001111101001: begin out_real=16'b0000001001000010; out_imag=16'b0011111111110110; end // in_theta = 0.488770 pi
 12'b001111101010: begin out_real=16'b0000001000101001; out_imag=16'b0011111111110111; end // in_theta = 0.489258 pi
 12'b001111101011: begin out_real=16'b0000001000010000; out_imag=16'b0011111111110111; end // in_theta = 0.489746 pi
 12'b001111101100: begin out_real=16'b0000000111110111; out_imag=16'b0011111111111000; end // in_theta = 0.490234 pi
 12'b001111101101: begin out_real=16'b0000000111011101; out_imag=16'b0011111111111001; end // in_theta = 0.490723 pi
 12'b001111101110: begin out_real=16'b0000000111000100; out_imag=16'b0011111111111010; end // in_theta = 0.491211 pi
 12'b001111101111: begin out_real=16'b0000000110101011; out_imag=16'b0011111111111010; end // in_theta = 0.491699 pi
 12'b001111110000: begin out_real=16'b0000000110010010; out_imag=16'b0011111111111011; end // in_theta = 0.492188 pi
 12'b001111110001: begin out_real=16'b0000000101111001; out_imag=16'b0011111111111100; end // in_theta = 0.492676 pi
 12'b001111110010: begin out_real=16'b0000000101100000; out_imag=16'b0011111111111100; end // in_theta = 0.493164 pi
 12'b001111110011: begin out_real=16'b0000000101000111; out_imag=16'b0011111111111101; end // in_theta = 0.493652 pi
 12'b001111110100: begin out_real=16'b0000000100101110; out_imag=16'b0011111111111101; end // in_theta = 0.494141 pi
 12'b001111110101: begin out_real=16'b0000000100010100; out_imag=16'b0011111111111110; end // in_theta = 0.494629 pi
 12'b001111110110: begin out_real=16'b0000000011111011; out_imag=16'b0011111111111110; end // in_theta = 0.495117 pi
 12'b001111110111: begin out_real=16'b0000000011100010; out_imag=16'b0011111111111110; end // in_theta = 0.495605 pi
 12'b001111111000: begin out_real=16'b0000000011001001; out_imag=16'b0011111111111111; end // in_theta = 0.496094 pi
 12'b001111111001: begin out_real=16'b0000000010110000; out_imag=16'b0011111111111111; end // in_theta = 0.496582 pi
 12'b001111111010: begin out_real=16'b0000000010010111; out_imag=16'b0011111111111111; end // in_theta = 0.497070 pi
 12'b001111111011: begin out_real=16'b0000000001111110; out_imag=16'b0100000000000000; end // in_theta = 0.497559 pi
 12'b001111111100: begin out_real=16'b0000000001100101; out_imag=16'b0100000000000000; end // in_theta = 0.498047 pi
 12'b001111111101: begin out_real=16'b0000000001001011; out_imag=16'b0100000000000000; end // in_theta = 0.498535 pi
 12'b001111111110: begin out_real=16'b0000000000110010; out_imag=16'b0100000000000000; end // in_theta = 0.499023 pi
 12'b001111111111: begin out_real=16'b0000000000011001; out_imag=16'b0100000000000000; end // in_theta = 0.499512 pi
 12'b010000000000: begin out_real=16'b0000000000000000; out_imag=16'b0100000000000000; end // in_theta = 0.500000 pi
 12'b010000000001: begin out_real=16'b1111111111100111; out_imag=16'b0100000000000000; end // in_theta = 0.500488 pi
 12'b010000000010: begin out_real=16'b1111111111001110; out_imag=16'b0100000000000000; end // in_theta = 0.500977 pi
 12'b010000000011: begin out_real=16'b1111111110110101; out_imag=16'b0100000000000000; end // in_theta = 0.501465 pi
 12'b010000000100: begin out_real=16'b1111111110011011; out_imag=16'b0100000000000000; end // in_theta = 0.501953 pi
 12'b010000000101: begin out_real=16'b1111111110000010; out_imag=16'b0100000000000000; end // in_theta = 0.502441 pi
 12'b010000000110: begin out_real=16'b1111111101101001; out_imag=16'b0011111111111111; end // in_theta = 0.502930 pi
 12'b010000000111: begin out_real=16'b1111111101010000; out_imag=16'b0011111111111111; end // in_theta = 0.503418 pi
 12'b010000001000: begin out_real=16'b1111111100110111; out_imag=16'b0011111111111111; end // in_theta = 0.503906 pi
 12'b010000001001: begin out_real=16'b1111111100011110; out_imag=16'b0011111111111110; end // in_theta = 0.504395 pi
 12'b010000001010: begin out_real=16'b1111111100000101; out_imag=16'b0011111111111110; end // in_theta = 0.504883 pi
 12'b010000001011: begin out_real=16'b1111111011101100; out_imag=16'b0011111111111110; end // in_theta = 0.505371 pi
 12'b010000001100: begin out_real=16'b1111111011010010; out_imag=16'b0011111111111101; end // in_theta = 0.505859 pi
 12'b010000001101: begin out_real=16'b1111111010111001; out_imag=16'b0011111111111101; end // in_theta = 0.506348 pi
 12'b010000001110: begin out_real=16'b1111111010100000; out_imag=16'b0011111111111100; end // in_theta = 0.506836 pi
 12'b010000001111: begin out_real=16'b1111111010000111; out_imag=16'b0011111111111100; end // in_theta = 0.507324 pi
 12'b010000010000: begin out_real=16'b1111111001101110; out_imag=16'b0011111111111011; end // in_theta = 0.507813 pi
 12'b010000010001: begin out_real=16'b1111111001010101; out_imag=16'b0011111111111010; end // in_theta = 0.508301 pi
 12'b010000010010: begin out_real=16'b1111111000111100; out_imag=16'b0011111111111010; end // in_theta = 0.508789 pi
 12'b010000010011: begin out_real=16'b1111111000100011; out_imag=16'b0011111111111001; end // in_theta = 0.509277 pi
 12'b010000010100: begin out_real=16'b1111111000001001; out_imag=16'b0011111111111000; end // in_theta = 0.509766 pi
 12'b010000010101: begin out_real=16'b1111110111110000; out_imag=16'b0011111111110111; end // in_theta = 0.510254 pi
 12'b010000010110: begin out_real=16'b1111110111010111; out_imag=16'b0011111111110111; end // in_theta = 0.510742 pi
 12'b010000010111: begin out_real=16'b1111110110111110; out_imag=16'b0011111111110110; end // in_theta = 0.511230 pi
 12'b010000011000: begin out_real=16'b1111110110100101; out_imag=16'b0011111111110101; end // in_theta = 0.511719 pi
 12'b010000011001: begin out_real=16'b1111110110001100; out_imag=16'b0011111111110100; end // in_theta = 0.512207 pi
 12'b010000011010: begin out_real=16'b1111110101110011; out_imag=16'b0011111111110011; end // in_theta = 0.512695 pi
 12'b010000011011: begin out_real=16'b1111110101011010; out_imag=16'b0011111111110010; end // in_theta = 0.513184 pi
 12'b010000011100: begin out_real=16'b1111110101000000; out_imag=16'b0011111111110001; end // in_theta = 0.513672 pi
 12'b010000011101: begin out_real=16'b1111110100100111; out_imag=16'b0011111111110000; end // in_theta = 0.514160 pi
 12'b010000011110: begin out_real=16'b1111110100001110; out_imag=16'b0011111111101111; end // in_theta = 0.514648 pi
 12'b010000011111: begin out_real=16'b1111110011110101; out_imag=16'b0011111111101101; end // in_theta = 0.515137 pi
 12'b010000100000: begin out_real=16'b1111110011011100; out_imag=16'b0011111111101100; end // in_theta = 0.515625 pi
 12'b010000100001: begin out_real=16'b1111110011000011; out_imag=16'b0011111111101011; end // in_theta = 0.516113 pi
 12'b010000100010: begin out_real=16'b1111110010101010; out_imag=16'b0011111111101010; end // in_theta = 0.516602 pi
 12'b010000100011: begin out_real=16'b1111110010010001; out_imag=16'b0011111111101000; end // in_theta = 0.517090 pi
 12'b010000100100: begin out_real=16'b1111110001111000; out_imag=16'b0011111111100111; end // in_theta = 0.517578 pi
 12'b010000100101: begin out_real=16'b1111110001011111; out_imag=16'b0011111111100110; end // in_theta = 0.518066 pi
 12'b010000100110: begin out_real=16'b1111110001000101; out_imag=16'b0011111111100100; end // in_theta = 0.518555 pi
 12'b010000100111: begin out_real=16'b1111110000101100; out_imag=16'b0011111111100011; end // in_theta = 0.519043 pi
 12'b010000101000: begin out_real=16'b1111110000010011; out_imag=16'b0011111111100001; end // in_theta = 0.519531 pi
 12'b010000101001: begin out_real=16'b1111101111111010; out_imag=16'b0011111111100000; end // in_theta = 0.520020 pi
 12'b010000101010: begin out_real=16'b1111101111100001; out_imag=16'b0011111111011110; end // in_theta = 0.520508 pi
 12'b010000101011: begin out_real=16'b1111101111001000; out_imag=16'b0011111111011100; end // in_theta = 0.520996 pi
 12'b010000101100: begin out_real=16'b1111101110101111; out_imag=16'b0011111111011011; end // in_theta = 0.521484 pi
 12'b010000101101: begin out_real=16'b1111101110010110; out_imag=16'b0011111111011001; end // in_theta = 0.521973 pi
 12'b010000101110: begin out_real=16'b1111101101111101; out_imag=16'b0011111111010111; end // in_theta = 0.522461 pi
 12'b010000101111: begin out_real=16'b1111101101100100; out_imag=16'b0011111111010101; end // in_theta = 0.522949 pi
 12'b010000110000: begin out_real=16'b1111101101001011; out_imag=16'b0011111111010100; end // in_theta = 0.523438 pi
 12'b010000110001: begin out_real=16'b1111101100110010; out_imag=16'b0011111111010010; end // in_theta = 0.523926 pi
 12'b010000110010: begin out_real=16'b1111101100011001; out_imag=16'b0011111111010000; end // in_theta = 0.524414 pi
 12'b010000110011: begin out_real=16'b1111101100000000; out_imag=16'b0011111111001110; end // in_theta = 0.524902 pi
 12'b010000110100: begin out_real=16'b1111101011100110; out_imag=16'b0011111111001100; end // in_theta = 0.525391 pi
 12'b010000110101: begin out_real=16'b1111101011001101; out_imag=16'b0011111111001010; end // in_theta = 0.525879 pi
 12'b010000110110: begin out_real=16'b1111101010110100; out_imag=16'b0011111111001000; end // in_theta = 0.526367 pi
 12'b010000110111: begin out_real=16'b1111101010011011; out_imag=16'b0011111111000110; end // in_theta = 0.526855 pi
 12'b010000111000: begin out_real=16'b1111101010000010; out_imag=16'b0011111111000100; end // in_theta = 0.527344 pi
 12'b010000111001: begin out_real=16'b1111101001101001; out_imag=16'b0011111111000001; end // in_theta = 0.527832 pi
 12'b010000111010: begin out_real=16'b1111101001010000; out_imag=16'b0011111110111111; end // in_theta = 0.528320 pi
 12'b010000111011: begin out_real=16'b1111101000110111; out_imag=16'b0011111110111101; end // in_theta = 0.528809 pi
 12'b010000111100: begin out_real=16'b1111101000011110; out_imag=16'b0011111110111011; end // in_theta = 0.529297 pi
 12'b010000111101: begin out_real=16'b1111101000000101; out_imag=16'b0011111110111000; end // in_theta = 0.529785 pi
 12'b010000111110: begin out_real=16'b1111100111101100; out_imag=16'b0011111110110110; end // in_theta = 0.530273 pi
 12'b010000111111: begin out_real=16'b1111100111010011; out_imag=16'b0011111110110100; end // in_theta = 0.530762 pi
 12'b010001000000: begin out_real=16'b1111100110111010; out_imag=16'b0011111110110001; end // in_theta = 0.531250 pi
 12'b010001000001: begin out_real=16'b1111100110100001; out_imag=16'b0011111110101111; end // in_theta = 0.531738 pi
 12'b010001000010: begin out_real=16'b1111100110001000; out_imag=16'b0011111110101100; end // in_theta = 0.532227 pi
 12'b010001000011: begin out_real=16'b1111100101101111; out_imag=16'b0011111110101010; end // in_theta = 0.532715 pi
 12'b010001000100: begin out_real=16'b1111100101010110; out_imag=16'b0011111110100111; end // in_theta = 0.533203 pi
 12'b010001000101: begin out_real=16'b1111100100111101; out_imag=16'b0011111110100100; end // in_theta = 0.533691 pi
 12'b010001000110: begin out_real=16'b1111100100100100; out_imag=16'b0011111110100010; end // in_theta = 0.534180 pi
 12'b010001000111: begin out_real=16'b1111100100001011; out_imag=16'b0011111110011111; end // in_theta = 0.534668 pi
 12'b010001001000: begin out_real=16'b1111100011110010; out_imag=16'b0011111110011100; end // in_theta = 0.535156 pi
 12'b010001001001: begin out_real=16'b1111100011011001; out_imag=16'b0011111110011001; end // in_theta = 0.535645 pi
 12'b010001001010: begin out_real=16'b1111100011000000; out_imag=16'b0011111110010111; end // in_theta = 0.536133 pi
 12'b010001001011: begin out_real=16'b1111100010100111; out_imag=16'b0011111110010100; end // in_theta = 0.536621 pi
 12'b010001001100: begin out_real=16'b1111100010001110; out_imag=16'b0011111110010001; end // in_theta = 0.537109 pi
 12'b010001001101: begin out_real=16'b1111100001110101; out_imag=16'b0011111110001110; end // in_theta = 0.537598 pi
 12'b010001001110: begin out_real=16'b1111100001011100; out_imag=16'b0011111110001011; end // in_theta = 0.538086 pi
 12'b010001001111: begin out_real=16'b1111100001000011; out_imag=16'b0011111110001000; end // in_theta = 0.538574 pi
 12'b010001010000: begin out_real=16'b1111100000101010; out_imag=16'b0011111110000101; end // in_theta = 0.539063 pi
 12'b010001010001: begin out_real=16'b1111100000010001; out_imag=16'b0011111110000010; end // in_theta = 0.539551 pi
 12'b010001010010: begin out_real=16'b1111011111111001; out_imag=16'b0011111101111111; end // in_theta = 0.540039 pi
 12'b010001010011: begin out_real=16'b1111011111100000; out_imag=16'b0011111101111011; end // in_theta = 0.540527 pi
 12'b010001010100: begin out_real=16'b1111011111000111; out_imag=16'b0011111101111000; end // in_theta = 0.541016 pi
 12'b010001010101: begin out_real=16'b1111011110101110; out_imag=16'b0011111101110101; end // in_theta = 0.541504 pi
 12'b010001010110: begin out_real=16'b1111011110010101; out_imag=16'b0011111101110010; end // in_theta = 0.541992 pi
 12'b010001010111: begin out_real=16'b1111011101111100; out_imag=16'b0011111101101110; end // in_theta = 0.542480 pi
 12'b010001011000: begin out_real=16'b1111011101100011; out_imag=16'b0011111101101011; end // in_theta = 0.542969 pi
 12'b010001011001: begin out_real=16'b1111011101001010; out_imag=16'b0011111101101000; end // in_theta = 0.543457 pi
 12'b010001011010: begin out_real=16'b1111011100110001; out_imag=16'b0011111101100100; end // in_theta = 0.543945 pi
 12'b010001011011: begin out_real=16'b1111011100011000; out_imag=16'b0011111101100001; end // in_theta = 0.544434 pi
 12'b010001011100: begin out_real=16'b1111011011111111; out_imag=16'b0011111101011101; end // in_theta = 0.544922 pi
 12'b010001011101: begin out_real=16'b1111011011100111; out_imag=16'b0011111101011010; end // in_theta = 0.545410 pi
 12'b010001011110: begin out_real=16'b1111011011001110; out_imag=16'b0011111101010110; end // in_theta = 0.545898 pi
 12'b010001011111: begin out_real=16'b1111011010110101; out_imag=16'b0011111101010010; end // in_theta = 0.546387 pi
 12'b010001100000: begin out_real=16'b1111011010011100; out_imag=16'b0011111101001111; end // in_theta = 0.546875 pi
 12'b010001100001: begin out_real=16'b1111011010000011; out_imag=16'b0011111101001011; end // in_theta = 0.547363 pi
 12'b010001100010: begin out_real=16'b1111011001101010; out_imag=16'b0011111101000111; end // in_theta = 0.547852 pi
 12'b010001100011: begin out_real=16'b1111011001010001; out_imag=16'b0011111101000011; end // in_theta = 0.548340 pi
 12'b010001100100: begin out_real=16'b1111011000111001; out_imag=16'b0011111101000000; end // in_theta = 0.548828 pi
 12'b010001100101: begin out_real=16'b1111011000100000; out_imag=16'b0011111100111100; end // in_theta = 0.549316 pi
 12'b010001100110: begin out_real=16'b1111011000000111; out_imag=16'b0011111100111000; end // in_theta = 0.549805 pi
 12'b010001100111: begin out_real=16'b1111010111101110; out_imag=16'b0011111100110100; end // in_theta = 0.550293 pi
 12'b010001101000: begin out_real=16'b1111010111010101; out_imag=16'b0011111100110000; end // in_theta = 0.550781 pi
 12'b010001101001: begin out_real=16'b1111010110111100; out_imag=16'b0011111100101100; end // in_theta = 0.551270 pi
 12'b010001101010: begin out_real=16'b1111010110100100; out_imag=16'b0011111100101000; end // in_theta = 0.551758 pi
 12'b010001101011: begin out_real=16'b1111010110001011; out_imag=16'b0011111100100100; end // in_theta = 0.552246 pi
 12'b010001101100: begin out_real=16'b1111010101110010; out_imag=16'b0011111100100000; end // in_theta = 0.552734 pi
 12'b010001101101: begin out_real=16'b1111010101011001; out_imag=16'b0011111100011100; end // in_theta = 0.553223 pi
 12'b010001101110: begin out_real=16'b1111010101000000; out_imag=16'b0011111100010111; end // in_theta = 0.553711 pi
 12'b010001101111: begin out_real=16'b1111010100101000; out_imag=16'b0011111100010011; end // in_theta = 0.554199 pi
 12'b010001110000: begin out_real=16'b1111010100001111; out_imag=16'b0011111100001111; end // in_theta = 0.554688 pi
 12'b010001110001: begin out_real=16'b1111010011110110; out_imag=16'b0011111100001010; end // in_theta = 0.555176 pi
 12'b010001110010: begin out_real=16'b1111010011011101; out_imag=16'b0011111100000110; end // in_theta = 0.555664 pi
 12'b010001110011: begin out_real=16'b1111010011000101; out_imag=16'b0011111100000010; end // in_theta = 0.556152 pi
 12'b010001110100: begin out_real=16'b1111010010101100; out_imag=16'b0011111011111101; end // in_theta = 0.556641 pi
 12'b010001110101: begin out_real=16'b1111010010010011; out_imag=16'b0011111011111001; end // in_theta = 0.557129 pi
 12'b010001110110: begin out_real=16'b1111010001111011; out_imag=16'b0011111011110100; end // in_theta = 0.557617 pi
 12'b010001110111: begin out_real=16'b1111010001100010; out_imag=16'b0011111011110000; end // in_theta = 0.558105 pi
 12'b010001111000: begin out_real=16'b1111010001001001; out_imag=16'b0011111011101011; end // in_theta = 0.558594 pi
 12'b010001111001: begin out_real=16'b1111010000110000; out_imag=16'b0011111011100111; end // in_theta = 0.559082 pi
 12'b010001111010: begin out_real=16'b1111010000011000; out_imag=16'b0011111011100010; end // in_theta = 0.559570 pi
 12'b010001111011: begin out_real=16'b1111001111111111; out_imag=16'b0011111011011101; end // in_theta = 0.560059 pi
 12'b010001111100: begin out_real=16'b1111001111100110; out_imag=16'b0011111011011000; end // in_theta = 0.560547 pi
 12'b010001111101: begin out_real=16'b1111001111001110; out_imag=16'b0011111011010100; end // in_theta = 0.561035 pi
 12'b010001111110: begin out_real=16'b1111001110110101; out_imag=16'b0011111011001111; end // in_theta = 0.561523 pi
 12'b010001111111: begin out_real=16'b1111001110011100; out_imag=16'b0011111011001010; end // in_theta = 0.562012 pi
 12'b010010000000: begin out_real=16'b1111001110000100; out_imag=16'b0011111011000101; end // in_theta = 0.562500 pi
 12'b010010000001: begin out_real=16'b1111001101101011; out_imag=16'b0011111011000000; end // in_theta = 0.562988 pi
 12'b010010000010: begin out_real=16'b1111001101010010; out_imag=16'b0011111010111011; end // in_theta = 0.563477 pi
 12'b010010000011: begin out_real=16'b1111001100111010; out_imag=16'b0011111010110110; end // in_theta = 0.563965 pi
 12'b010010000100: begin out_real=16'b1111001100100001; out_imag=16'b0011111010110001; end // in_theta = 0.564453 pi
 12'b010010000101: begin out_real=16'b1111001100001000; out_imag=16'b0011111010101100; end // in_theta = 0.564941 pi
 12'b010010000110: begin out_real=16'b1111001011110000; out_imag=16'b0011111010100111; end // in_theta = 0.565430 pi
 12'b010010000111: begin out_real=16'b1111001011010111; out_imag=16'b0011111010100010; end // in_theta = 0.565918 pi
 12'b010010001000: begin out_real=16'b1111001010111111; out_imag=16'b0011111010011101; end // in_theta = 0.566406 pi
 12'b010010001001: begin out_real=16'b1111001010100110; out_imag=16'b0011111010011000; end // in_theta = 0.566895 pi
 12'b010010001010: begin out_real=16'b1111001010001110; out_imag=16'b0011111010010010; end // in_theta = 0.567383 pi
 12'b010010001011: begin out_real=16'b1111001001110101; out_imag=16'b0011111010001101; end // in_theta = 0.567871 pi
 12'b010010001100: begin out_real=16'b1111001001011100; out_imag=16'b0011111010001000; end // in_theta = 0.568359 pi
 12'b010010001101: begin out_real=16'b1111001001000100; out_imag=16'b0011111010000010; end // in_theta = 0.568848 pi
 12'b010010001110: begin out_real=16'b1111001000101011; out_imag=16'b0011111001111101; end // in_theta = 0.569336 pi
 12'b010010001111: begin out_real=16'b1111001000010011; out_imag=16'b0011111001110111; end // in_theta = 0.569824 pi
 12'b010010010000: begin out_real=16'b1111000111111010; out_imag=16'b0011111001110010; end // in_theta = 0.570313 pi
 12'b010010010001: begin out_real=16'b1111000111100010; out_imag=16'b0011111001101100; end // in_theta = 0.570801 pi
 12'b010010010010: begin out_real=16'b1111000111001001; out_imag=16'b0011111001100111; end // in_theta = 0.571289 pi
 12'b010010010011: begin out_real=16'b1111000110110001; out_imag=16'b0011111001100001; end // in_theta = 0.571777 pi
 12'b010010010100: begin out_real=16'b1111000110011000; out_imag=16'b0011111001011100; end // in_theta = 0.572266 pi
 12'b010010010101: begin out_real=16'b1111000110000000; out_imag=16'b0011111001010110; end // in_theta = 0.572754 pi
 12'b010010010110: begin out_real=16'b1111000101100111; out_imag=16'b0011111001010000; end // in_theta = 0.573242 pi
 12'b010010010111: begin out_real=16'b1111000101001111; out_imag=16'b0011111001001010; end // in_theta = 0.573730 pi
 12'b010010011000: begin out_real=16'b1111000100110110; out_imag=16'b0011111001000101; end // in_theta = 0.574219 pi
 12'b010010011001: begin out_real=16'b1111000100011110; out_imag=16'b0011111000111111; end // in_theta = 0.574707 pi
 12'b010010011010: begin out_real=16'b1111000100000101; out_imag=16'b0011111000111001; end // in_theta = 0.575195 pi
 12'b010010011011: begin out_real=16'b1111000011101101; out_imag=16'b0011111000110011; end // in_theta = 0.575684 pi
 12'b010010011100: begin out_real=16'b1111000011010101; out_imag=16'b0011111000101101; end // in_theta = 0.576172 pi
 12'b010010011101: begin out_real=16'b1111000010111100; out_imag=16'b0011111000100111; end // in_theta = 0.576660 pi
 12'b010010011110: begin out_real=16'b1111000010100100; out_imag=16'b0011111000100001; end // in_theta = 0.577148 pi
 12'b010010011111: begin out_real=16'b1111000010001011; out_imag=16'b0011111000011011; end // in_theta = 0.577637 pi
 12'b010010100000: begin out_real=16'b1111000001110011; out_imag=16'b0011111000010101; end // in_theta = 0.578125 pi
 12'b010010100001: begin out_real=16'b1111000001011011; out_imag=16'b0011111000001111; end // in_theta = 0.578613 pi
 12'b010010100010: begin out_real=16'b1111000001000010; out_imag=16'b0011111000001001; end // in_theta = 0.579102 pi
 12'b010010100011: begin out_real=16'b1111000000101010; out_imag=16'b0011111000000011; end // in_theta = 0.579590 pi
 12'b010010100100: begin out_real=16'b1111000000010010; out_imag=16'b0011110111111100; end // in_theta = 0.580078 pi
 12'b010010100101: begin out_real=16'b1110111111111001; out_imag=16'b0011110111110110; end // in_theta = 0.580566 pi
 12'b010010100110: begin out_real=16'b1110111111100001; out_imag=16'b0011110111110000; end // in_theta = 0.581055 pi
 12'b010010100111: begin out_real=16'b1110111111001001; out_imag=16'b0011110111101001; end // in_theta = 0.581543 pi
 12'b010010101000: begin out_real=16'b1110111110110000; out_imag=16'b0011110111100011; end // in_theta = 0.582031 pi
 12'b010010101001: begin out_real=16'b1110111110011000; out_imag=16'b0011110111011101; end // in_theta = 0.582520 pi
 12'b010010101010: begin out_real=16'b1110111110000000; out_imag=16'b0011110111010110; end // in_theta = 0.583008 pi
 12'b010010101011: begin out_real=16'b1110111101100111; out_imag=16'b0011110111010000; end // in_theta = 0.583496 pi
 12'b010010101100: begin out_real=16'b1110111101001111; out_imag=16'b0011110111001001; end // in_theta = 0.583984 pi
 12'b010010101101: begin out_real=16'b1110111100110111; out_imag=16'b0011110111000010; end // in_theta = 0.584473 pi
 12'b010010101110: begin out_real=16'b1110111100011111; out_imag=16'b0011110110111100; end // in_theta = 0.584961 pi
 12'b010010101111: begin out_real=16'b1110111100000110; out_imag=16'b0011110110110101; end // in_theta = 0.585449 pi
 12'b010010110000: begin out_real=16'b1110111011101110; out_imag=16'b0011110110101111; end // in_theta = 0.585938 pi
 12'b010010110001: begin out_real=16'b1110111011010110; out_imag=16'b0011110110101000; end // in_theta = 0.586426 pi
 12'b010010110010: begin out_real=16'b1110111010111110; out_imag=16'b0011110110100001; end // in_theta = 0.586914 pi
 12'b010010110011: begin out_real=16'b1110111010100110; out_imag=16'b0011110110011010; end // in_theta = 0.587402 pi
 12'b010010110100: begin out_real=16'b1110111010001101; out_imag=16'b0011110110010011; end // in_theta = 0.587891 pi
 12'b010010110101: begin out_real=16'b1110111001110101; out_imag=16'b0011110110001101; end // in_theta = 0.588379 pi
 12'b010010110110: begin out_real=16'b1110111001011101; out_imag=16'b0011110110000110; end // in_theta = 0.588867 pi
 12'b010010110111: begin out_real=16'b1110111001000101; out_imag=16'b0011110101111111; end // in_theta = 0.589355 pi
 12'b010010111000: begin out_real=16'b1110111000101101; out_imag=16'b0011110101111000; end // in_theta = 0.589844 pi
 12'b010010111001: begin out_real=16'b1110111000010101; out_imag=16'b0011110101110001; end // in_theta = 0.590332 pi
 12'b010010111010: begin out_real=16'b1110110111111100; out_imag=16'b0011110101101010; end // in_theta = 0.590820 pi
 12'b010010111011: begin out_real=16'b1110110111100100; out_imag=16'b0011110101100011; end // in_theta = 0.591309 pi
 12'b010010111100: begin out_real=16'b1110110111001100; out_imag=16'b0011110101011011; end // in_theta = 0.591797 pi
 12'b010010111101: begin out_real=16'b1110110110110100; out_imag=16'b0011110101010100; end // in_theta = 0.592285 pi
 12'b010010111110: begin out_real=16'b1110110110011100; out_imag=16'b0011110101001101; end // in_theta = 0.592773 pi
 12'b010010111111: begin out_real=16'b1110110110000100; out_imag=16'b0011110101000110; end // in_theta = 0.593262 pi
 12'b010011000000: begin out_real=16'b1110110101101100; out_imag=16'b0011110100111111; end // in_theta = 0.593750 pi
 12'b010011000001: begin out_real=16'b1110110101010100; out_imag=16'b0011110100110111; end // in_theta = 0.594238 pi
 12'b010011000010: begin out_real=16'b1110110100111100; out_imag=16'b0011110100110000; end // in_theta = 0.594727 pi
 12'b010011000011: begin out_real=16'b1110110100100100; out_imag=16'b0011110100101000; end // in_theta = 0.595215 pi
 12'b010011000100: begin out_real=16'b1110110100001100; out_imag=16'b0011110100100001; end // in_theta = 0.595703 pi
 12'b010011000101: begin out_real=16'b1110110011110100; out_imag=16'b0011110100011010; end // in_theta = 0.596191 pi
 12'b010011000110: begin out_real=16'b1110110011011100; out_imag=16'b0011110100010010; end // in_theta = 0.596680 pi
 12'b010011000111: begin out_real=16'b1110110011000100; out_imag=16'b0011110100001011; end // in_theta = 0.597168 pi
 12'b010011001000: begin out_real=16'b1110110010101100; out_imag=16'b0011110100000011; end // in_theta = 0.597656 pi
 12'b010011001001: begin out_real=16'b1110110010010100; out_imag=16'b0011110011111011; end // in_theta = 0.598145 pi
 12'b010011001010: begin out_real=16'b1110110001111100; out_imag=16'b0011110011110100; end // in_theta = 0.598633 pi
 12'b010011001011: begin out_real=16'b1110110001100100; out_imag=16'b0011110011101100; end // in_theta = 0.599121 pi
 12'b010011001100: begin out_real=16'b1110110001001100; out_imag=16'b0011110011100100; end // in_theta = 0.599609 pi
 12'b010011001101: begin out_real=16'b1110110000110100; out_imag=16'b0011110011011101; end // in_theta = 0.600098 pi
 12'b010011001110: begin out_real=16'b1110110000011100; out_imag=16'b0011110011010101; end // in_theta = 0.600586 pi
 12'b010011001111: begin out_real=16'b1110110000000101; out_imag=16'b0011110011001101; end // in_theta = 0.601074 pi
 12'b010011010000: begin out_real=16'b1110101111101101; out_imag=16'b0011110011000101; end // in_theta = 0.601563 pi
 12'b010011010001: begin out_real=16'b1110101111010101; out_imag=16'b0011110010111101; end // in_theta = 0.602051 pi
 12'b010011010010: begin out_real=16'b1110101110111101; out_imag=16'b0011110010110101; end // in_theta = 0.602539 pi
 12'b010011010011: begin out_real=16'b1110101110100101; out_imag=16'b0011110010101101; end // in_theta = 0.603027 pi
 12'b010011010100: begin out_real=16'b1110101110001101; out_imag=16'b0011110010100101; end // in_theta = 0.603516 pi
 12'b010011010101: begin out_real=16'b1110101101110101; out_imag=16'b0011110010011101; end // in_theta = 0.604004 pi
 12'b010011010110: begin out_real=16'b1110101101011110; out_imag=16'b0011110010010101; end // in_theta = 0.604492 pi
 12'b010011010111: begin out_real=16'b1110101101000110; out_imag=16'b0011110010001101; end // in_theta = 0.604980 pi
 12'b010011011000: begin out_real=16'b1110101100101110; out_imag=16'b0011110010000101; end // in_theta = 0.605469 pi
 12'b010011011001: begin out_real=16'b1110101100010110; out_imag=16'b0011110001111101; end // in_theta = 0.605957 pi
 12'b010011011010: begin out_real=16'b1110101011111111; out_imag=16'b0011110001110100; end // in_theta = 0.606445 pi
 12'b010011011011: begin out_real=16'b1110101011100111; out_imag=16'b0011110001101100; end // in_theta = 0.606934 pi
 12'b010011011100: begin out_real=16'b1110101011001111; out_imag=16'b0011110001100100; end // in_theta = 0.607422 pi
 12'b010011011101: begin out_real=16'b1110101010110111; out_imag=16'b0011110001011011; end // in_theta = 0.607910 pi
 12'b010011011110: begin out_real=16'b1110101010100000; out_imag=16'b0011110001010011; end // in_theta = 0.608398 pi
 12'b010011011111: begin out_real=16'b1110101010001000; out_imag=16'b0011110001001011; end // in_theta = 0.608887 pi
 12'b010011100000: begin out_real=16'b1110101001110000; out_imag=16'b0011110001000010; end // in_theta = 0.609375 pi
 12'b010011100001: begin out_real=16'b1110101001011001; out_imag=16'b0011110000111010; end // in_theta = 0.609863 pi
 12'b010011100010: begin out_real=16'b1110101001000001; out_imag=16'b0011110000110001; end // in_theta = 0.610352 pi
 12'b010011100011: begin out_real=16'b1110101000101001; out_imag=16'b0011110000101001; end // in_theta = 0.610840 pi
 12'b010011100100: begin out_real=16'b1110101000010010; out_imag=16'b0011110000100000; end // in_theta = 0.611328 pi
 12'b010011100101: begin out_real=16'b1110100111111010; out_imag=16'b0011110000010111; end // in_theta = 0.611816 pi
 12'b010011100110: begin out_real=16'b1110100111100011; out_imag=16'b0011110000001111; end // in_theta = 0.612305 pi
 12'b010011100111: begin out_real=16'b1110100111001011; out_imag=16'b0011110000000110; end // in_theta = 0.612793 pi
 12'b010011101000: begin out_real=16'b1110100110110100; out_imag=16'b0011101111111101; end // in_theta = 0.613281 pi
 12'b010011101001: begin out_real=16'b1110100110011100; out_imag=16'b0011101111110101; end // in_theta = 0.613770 pi
 12'b010011101010: begin out_real=16'b1110100110000100; out_imag=16'b0011101111101100; end // in_theta = 0.614258 pi
 12'b010011101011: begin out_real=16'b1110100101101101; out_imag=16'b0011101111100011; end // in_theta = 0.614746 pi
 12'b010011101100: begin out_real=16'b1110100101010101; out_imag=16'b0011101111011010; end // in_theta = 0.615234 pi
 12'b010011101101: begin out_real=16'b1110100100111110; out_imag=16'b0011101111010001; end // in_theta = 0.615723 pi
 12'b010011101110: begin out_real=16'b1110100100100110; out_imag=16'b0011101111001000; end // in_theta = 0.616211 pi
 12'b010011101111: begin out_real=16'b1110100100001111; out_imag=16'b0011101110111111; end // in_theta = 0.616699 pi
 12'b010011110000: begin out_real=16'b1110100011110111; out_imag=16'b0011101110110110; end // in_theta = 0.617188 pi
 12'b010011110001: begin out_real=16'b1110100011100000; out_imag=16'b0011101110101101; end // in_theta = 0.617676 pi
 12'b010011110010: begin out_real=16'b1110100011001001; out_imag=16'b0011101110100100; end // in_theta = 0.618164 pi
 12'b010011110011: begin out_real=16'b1110100010110001; out_imag=16'b0011101110011011; end // in_theta = 0.618652 pi
 12'b010011110100: begin out_real=16'b1110100010011010; out_imag=16'b0011101110010010; end // in_theta = 0.619141 pi
 12'b010011110101: begin out_real=16'b1110100010000010; out_imag=16'b0011101110001000; end // in_theta = 0.619629 pi
 12'b010011110110: begin out_real=16'b1110100001101011; out_imag=16'b0011101101111111; end // in_theta = 0.620117 pi
 12'b010011110111: begin out_real=16'b1110100001010100; out_imag=16'b0011101101110110; end // in_theta = 0.620605 pi
 12'b010011111000: begin out_real=16'b1110100000111100; out_imag=16'b0011101101101101; end // in_theta = 0.621094 pi
 12'b010011111001: begin out_real=16'b1110100000100101; out_imag=16'b0011101101100011; end // in_theta = 0.621582 pi
 12'b010011111010: begin out_real=16'b1110100000001110; out_imag=16'b0011101101011010; end // in_theta = 0.622070 pi
 12'b010011111011: begin out_real=16'b1110011111110110; out_imag=16'b0011101101010000; end // in_theta = 0.622559 pi
 12'b010011111100: begin out_real=16'b1110011111011111; out_imag=16'b0011101101000111; end // in_theta = 0.623047 pi
 12'b010011111101: begin out_real=16'b1110011111001000; out_imag=16'b0011101100111110; end // in_theta = 0.623535 pi
 12'b010011111110: begin out_real=16'b1110011110110001; out_imag=16'b0011101100110100; end // in_theta = 0.624023 pi
 12'b010011111111: begin out_real=16'b1110011110011001; out_imag=16'b0011101100101010; end // in_theta = 0.624512 pi
 12'b010100000000: begin out_real=16'b1110011110000010; out_imag=16'b0011101100100001; end // in_theta = 0.625000 pi
 12'b010100000001: begin out_real=16'b1110011101101011; out_imag=16'b0011101100010111; end // in_theta = 0.625488 pi
 12'b010100000010: begin out_real=16'b1110011101010100; out_imag=16'b0011101100001110; end // in_theta = 0.625977 pi
 12'b010100000011: begin out_real=16'b1110011100111101; out_imag=16'b0011101100000100; end // in_theta = 0.626465 pi
 12'b010100000100: begin out_real=16'b1110011100100101; out_imag=16'b0011101011111010; end // in_theta = 0.626953 pi
 12'b010100000101: begin out_real=16'b1110011100001110; out_imag=16'b0011101011110000; end // in_theta = 0.627441 pi
 12'b010100000110: begin out_real=16'b1110011011110111; out_imag=16'b0011101011100110; end // in_theta = 0.627930 pi
 12'b010100000111: begin out_real=16'b1110011011100000; out_imag=16'b0011101011011101; end // in_theta = 0.628418 pi
 12'b010100001000: begin out_real=16'b1110011011001001; out_imag=16'b0011101011010011; end // in_theta = 0.628906 pi
 12'b010100001001: begin out_real=16'b1110011010110010; out_imag=16'b0011101011001001; end // in_theta = 0.629395 pi
 12'b010100001010: begin out_real=16'b1110011010011011; out_imag=16'b0011101010111111; end // in_theta = 0.629883 pi
 12'b010100001011: begin out_real=16'b1110011010000100; out_imag=16'b0011101010110101; end // in_theta = 0.630371 pi
 12'b010100001100: begin out_real=16'b1110011001101101; out_imag=16'b0011101010101011; end // in_theta = 0.630859 pi
 12'b010100001101: begin out_real=16'b1110011001010110; out_imag=16'b0011101010100001; end // in_theta = 0.631348 pi
 12'b010100001110: begin out_real=16'b1110011000111111; out_imag=16'b0011101010010111; end // in_theta = 0.631836 pi
 12'b010100001111: begin out_real=16'b1110011000101000; out_imag=16'b0011101010001101; end // in_theta = 0.632324 pi
 12'b010100010000: begin out_real=16'b1110011000010001; out_imag=16'b0011101010000010; end // in_theta = 0.632813 pi
 12'b010100010001: begin out_real=16'b1110010111111010; out_imag=16'b0011101001111000; end // in_theta = 0.633301 pi
 12'b010100010010: begin out_real=16'b1110010111100011; out_imag=16'b0011101001101110; end // in_theta = 0.633789 pi
 12'b010100010011: begin out_real=16'b1110010111001100; out_imag=16'b0011101001100100; end // in_theta = 0.634277 pi
 12'b010100010100: begin out_real=16'b1110010110110101; out_imag=16'b0011101001011001; end // in_theta = 0.634766 pi
 12'b010100010101: begin out_real=16'b1110010110011110; out_imag=16'b0011101001001111; end // in_theta = 0.635254 pi
 12'b010100010110: begin out_real=16'b1110010110000111; out_imag=16'b0011101001000101; end // in_theta = 0.635742 pi
 12'b010100010111: begin out_real=16'b1110010101110000; out_imag=16'b0011101000111010; end // in_theta = 0.636230 pi
 12'b010100011000: begin out_real=16'b1110010101011001; out_imag=16'b0011101000110000; end // in_theta = 0.636719 pi
 12'b010100011001: begin out_real=16'b1110010101000010; out_imag=16'b0011101000100101; end // in_theta = 0.637207 pi
 12'b010100011010: begin out_real=16'b1110010100101100; out_imag=16'b0011101000011011; end // in_theta = 0.637695 pi
 12'b010100011011: begin out_real=16'b1110010100010101; out_imag=16'b0011101000010000; end // in_theta = 0.638184 pi
 12'b010100011100: begin out_real=16'b1110010011111110; out_imag=16'b0011101000000110; end // in_theta = 0.638672 pi
 12'b010100011101: begin out_real=16'b1110010011100111; out_imag=16'b0011100111111011; end // in_theta = 0.639160 pi
 12'b010100011110: begin out_real=16'b1110010011010000; out_imag=16'b0011100111110000; end // in_theta = 0.639648 pi
 12'b010100011111: begin out_real=16'b1110010010111010; out_imag=16'b0011100111100110; end // in_theta = 0.640137 pi
 12'b010100100000: begin out_real=16'b1110010010100011; out_imag=16'b0011100111011011; end // in_theta = 0.640625 pi
 12'b010100100001: begin out_real=16'b1110010010001100; out_imag=16'b0011100111010000; end // in_theta = 0.641113 pi
 12'b010100100010: begin out_real=16'b1110010001110110; out_imag=16'b0011100111000101; end // in_theta = 0.641602 pi
 12'b010100100011: begin out_real=16'b1110010001011111; out_imag=16'b0011100110111011; end // in_theta = 0.642090 pi
 12'b010100100100: begin out_real=16'b1110010001001000; out_imag=16'b0011100110110000; end // in_theta = 0.642578 pi
 12'b010100100101: begin out_real=16'b1110010000110010; out_imag=16'b0011100110100101; end // in_theta = 0.643066 pi
 12'b010100100110: begin out_real=16'b1110010000011011; out_imag=16'b0011100110011010; end // in_theta = 0.643555 pi
 12'b010100100111: begin out_real=16'b1110010000000100; out_imag=16'b0011100110001111; end // in_theta = 0.644043 pi
 12'b010100101000: begin out_real=16'b1110001111101110; out_imag=16'b0011100110000100; end // in_theta = 0.644531 pi
 12'b010100101001: begin out_real=16'b1110001111010111; out_imag=16'b0011100101111001; end // in_theta = 0.645020 pi
 12'b010100101010: begin out_real=16'b1110001111000001; out_imag=16'b0011100101101110; end // in_theta = 0.645508 pi
 12'b010100101011: begin out_real=16'b1110001110101010; out_imag=16'b0011100101100011; end // in_theta = 0.645996 pi
 12'b010100101100: begin out_real=16'b1110001110010100; out_imag=16'b0011100101011000; end // in_theta = 0.646484 pi
 12'b010100101101: begin out_real=16'b1110001101111101; out_imag=16'b0011100101001100; end // in_theta = 0.646973 pi
 12'b010100101110: begin out_real=16'b1110001101100111; out_imag=16'b0011100101000001; end // in_theta = 0.647461 pi
 12'b010100101111: begin out_real=16'b1110001101010000; out_imag=16'b0011100100110110; end // in_theta = 0.647949 pi
 12'b010100110000: begin out_real=16'b1110001100111010; out_imag=16'b0011100100101011; end // in_theta = 0.648438 pi
 12'b010100110001: begin out_real=16'b1110001100100011; out_imag=16'b0011100100011111; end // in_theta = 0.648926 pi
 12'b010100110010: begin out_real=16'b1110001100001101; out_imag=16'b0011100100010100; end // in_theta = 0.649414 pi
 12'b010100110011: begin out_real=16'b1110001011110110; out_imag=16'b0011100100001001; end // in_theta = 0.649902 pi
 12'b010100110100: begin out_real=16'b1110001011100000; out_imag=16'b0011100011111101; end // in_theta = 0.650391 pi
 12'b010100110101: begin out_real=16'b1110001011001010; out_imag=16'b0011100011110010; end // in_theta = 0.650879 pi
 12'b010100110110: begin out_real=16'b1110001010110011; out_imag=16'b0011100011100110; end // in_theta = 0.651367 pi
 12'b010100110111: begin out_real=16'b1110001010011101; out_imag=16'b0011100011011011; end // in_theta = 0.651855 pi
 12'b010100111000: begin out_real=16'b1110001010000111; out_imag=16'b0011100011001111; end // in_theta = 0.652344 pi
 12'b010100111001: begin out_real=16'b1110001001110000; out_imag=16'b0011100011000011; end // in_theta = 0.652832 pi
 12'b010100111010: begin out_real=16'b1110001001011010; out_imag=16'b0011100010111000; end // in_theta = 0.653320 pi
 12'b010100111011: begin out_real=16'b1110001001000100; out_imag=16'b0011100010101100; end // in_theta = 0.653809 pi
 12'b010100111100: begin out_real=16'b1110001000101101; out_imag=16'b0011100010100001; end // in_theta = 0.654297 pi
 12'b010100111101: begin out_real=16'b1110001000010111; out_imag=16'b0011100010010101; end // in_theta = 0.654785 pi
 12'b010100111110: begin out_real=16'b1110001000000001; out_imag=16'b0011100010001001; end // in_theta = 0.655273 pi
 12'b010100111111: begin out_real=16'b1110000111101011; out_imag=16'b0011100001111101; end // in_theta = 0.655762 pi
 12'b010101000000: begin out_real=16'b1110000111010101; out_imag=16'b0011100001110001; end // in_theta = 0.656250 pi
 12'b010101000001: begin out_real=16'b1110000110111110; out_imag=16'b0011100001100110; end // in_theta = 0.656738 pi
 12'b010101000010: begin out_real=16'b1110000110101000; out_imag=16'b0011100001011010; end // in_theta = 0.657227 pi
 12'b010101000011: begin out_real=16'b1110000110010010; out_imag=16'b0011100001001110; end // in_theta = 0.657715 pi
 12'b010101000100: begin out_real=16'b1110000101111100; out_imag=16'b0011100001000010; end // in_theta = 0.658203 pi
 12'b010101000101: begin out_real=16'b1110000101100110; out_imag=16'b0011100000110110; end // in_theta = 0.658691 pi
 12'b010101000110: begin out_real=16'b1110000101010000; out_imag=16'b0011100000101010; end // in_theta = 0.659180 pi
 12'b010101000111: begin out_real=16'b1110000100111010; out_imag=16'b0011100000011110; end // in_theta = 0.659668 pi
 12'b010101001000: begin out_real=16'b1110000100100100; out_imag=16'b0011100000010010; end // in_theta = 0.660156 pi
 12'b010101001001: begin out_real=16'b1110000100001110; out_imag=16'b0011100000000101; end // in_theta = 0.660645 pi
 12'b010101001010: begin out_real=16'b1110000011111000; out_imag=16'b0011011111111001; end // in_theta = 0.661133 pi
 12'b010101001011: begin out_real=16'b1110000011100010; out_imag=16'b0011011111101101; end // in_theta = 0.661621 pi
 12'b010101001100: begin out_real=16'b1110000011001100; out_imag=16'b0011011111100001; end // in_theta = 0.662109 pi
 12'b010101001101: begin out_real=16'b1110000010110110; out_imag=16'b0011011111010101; end // in_theta = 0.662598 pi
 12'b010101001110: begin out_real=16'b1110000010100000; out_imag=16'b0011011111001000; end // in_theta = 0.663086 pi
 12'b010101001111: begin out_real=16'b1110000010001010; out_imag=16'b0011011110111100; end // in_theta = 0.663574 pi
 12'b010101010000: begin out_real=16'b1110000001110100; out_imag=16'b0011011110110000; end // in_theta = 0.664063 pi
 12'b010101010001: begin out_real=16'b1110000001011110; out_imag=16'b0011011110100011; end // in_theta = 0.664551 pi
 12'b010101010010: begin out_real=16'b1110000001001001; out_imag=16'b0011011110010111; end // in_theta = 0.665039 pi
 12'b010101010011: begin out_real=16'b1110000000110011; out_imag=16'b0011011110001010; end // in_theta = 0.665527 pi
 12'b010101010100: begin out_real=16'b1110000000011101; out_imag=16'b0011011101111110; end // in_theta = 0.666016 pi
 12'b010101010101: begin out_real=16'b1110000000000111; out_imag=16'b0011011101110001; end // in_theta = 0.666504 pi
 12'b010101010110: begin out_real=16'b1101111111110001; out_imag=16'b0011011101100101; end // in_theta = 0.666992 pi
 12'b010101010111: begin out_real=16'b1101111111011100; out_imag=16'b0011011101011000; end // in_theta = 0.667480 pi
 12'b010101011000: begin out_real=16'b1101111111000110; out_imag=16'b0011011101001011; end // in_theta = 0.667969 pi
 12'b010101011001: begin out_real=16'b1101111110110000; out_imag=16'b0011011100111111; end // in_theta = 0.668457 pi
 12'b010101011010: begin out_real=16'b1101111110011011; out_imag=16'b0011011100110010; end // in_theta = 0.668945 pi
 12'b010101011011: begin out_real=16'b1101111110000101; out_imag=16'b0011011100100101; end // in_theta = 0.669434 pi
 12'b010101011100: begin out_real=16'b1101111101101111; out_imag=16'b0011011100011000; end // in_theta = 0.669922 pi
 12'b010101011101: begin out_real=16'b1101111101011010; out_imag=16'b0011011100001100; end // in_theta = 0.670410 pi
 12'b010101011110: begin out_real=16'b1101111101000100; out_imag=16'b0011011011111111; end // in_theta = 0.670898 pi
 12'b010101011111: begin out_real=16'b1101111100101111; out_imag=16'b0011011011110010; end // in_theta = 0.671387 pi
 12'b010101100000: begin out_real=16'b1101111100011001; out_imag=16'b0011011011100101; end // in_theta = 0.671875 pi
 12'b010101100001: begin out_real=16'b1101111100000011; out_imag=16'b0011011011011000; end // in_theta = 0.672363 pi
 12'b010101100010: begin out_real=16'b1101111011101110; out_imag=16'b0011011011001011; end // in_theta = 0.672852 pi
 12'b010101100011: begin out_real=16'b1101111011011000; out_imag=16'b0011011010111110; end // in_theta = 0.673340 pi
 12'b010101100100: begin out_real=16'b1101111011000011; out_imag=16'b0011011010110001; end // in_theta = 0.673828 pi
 12'b010101100101: begin out_real=16'b1101111010101101; out_imag=16'b0011011010100100; end // in_theta = 0.674316 pi
 12'b010101100110: begin out_real=16'b1101111010011000; out_imag=16'b0011011010010111; end // in_theta = 0.674805 pi
 12'b010101100111: begin out_real=16'b1101111010000011; out_imag=16'b0011011010001010; end // in_theta = 0.675293 pi
 12'b010101101000: begin out_real=16'b1101111001101101; out_imag=16'b0011011001111101; end // in_theta = 0.675781 pi
 12'b010101101001: begin out_real=16'b1101111001011000; out_imag=16'b0011011001101111; end // in_theta = 0.676270 pi
 12'b010101101010: begin out_real=16'b1101111001000010; out_imag=16'b0011011001100010; end // in_theta = 0.676758 pi
 12'b010101101011: begin out_real=16'b1101111000101101; out_imag=16'b0011011001010101; end // in_theta = 0.677246 pi
 12'b010101101100: begin out_real=16'b1101111000011000; out_imag=16'b0011011001001000; end // in_theta = 0.677734 pi
 12'b010101101101: begin out_real=16'b1101111000000010; out_imag=16'b0011011000111010; end // in_theta = 0.678223 pi
 12'b010101101110: begin out_real=16'b1101110111101101; out_imag=16'b0011011000101101; end // in_theta = 0.678711 pi
 12'b010101101111: begin out_real=16'b1101110111011000; out_imag=16'b0011011000100000; end // in_theta = 0.679199 pi
 12'b010101110000: begin out_real=16'b1101110111000011; out_imag=16'b0011011000010010; end // in_theta = 0.679688 pi
 12'b010101110001: begin out_real=16'b1101110110101101; out_imag=16'b0011011000000101; end // in_theta = 0.680176 pi
 12'b010101110010: begin out_real=16'b1101110110011000; out_imag=16'b0011010111110111; end // in_theta = 0.680664 pi
 12'b010101110011: begin out_real=16'b1101110110000011; out_imag=16'b0011010111101010; end // in_theta = 0.681152 pi
 12'b010101110100: begin out_real=16'b1101110101101110; out_imag=16'b0011010111011100; end // in_theta = 0.681641 pi
 12'b010101110101: begin out_real=16'b1101110101011001; out_imag=16'b0011010111001110; end // in_theta = 0.682129 pi
 12'b010101110110: begin out_real=16'b1101110101000100; out_imag=16'b0011010111000001; end // in_theta = 0.682617 pi
 12'b010101110111: begin out_real=16'b1101110100101110; out_imag=16'b0011010110110011; end // in_theta = 0.683105 pi
 12'b010101111000: begin out_real=16'b1101110100011001; out_imag=16'b0011010110100101; end // in_theta = 0.683594 pi
 12'b010101111001: begin out_real=16'b1101110100000100; out_imag=16'b0011010110011000; end // in_theta = 0.684082 pi
 12'b010101111010: begin out_real=16'b1101110011101111; out_imag=16'b0011010110001010; end // in_theta = 0.684570 pi
 12'b010101111011: begin out_real=16'b1101110011011010; out_imag=16'b0011010101111100; end // in_theta = 0.685059 pi
 12'b010101111100: begin out_real=16'b1101110011000101; out_imag=16'b0011010101101110; end // in_theta = 0.685547 pi
 12'b010101111101: begin out_real=16'b1101110010110000; out_imag=16'b0011010101100001; end // in_theta = 0.686035 pi
 12'b010101111110: begin out_real=16'b1101110010011011; out_imag=16'b0011010101010011; end // in_theta = 0.686523 pi
 12'b010101111111: begin out_real=16'b1101110010000110; out_imag=16'b0011010101000101; end // in_theta = 0.687012 pi
 12'b010110000000: begin out_real=16'b1101110001110010; out_imag=16'b0011010100110111; end // in_theta = 0.687500 pi
 12'b010110000001: begin out_real=16'b1101110001011101; out_imag=16'b0011010100101001; end // in_theta = 0.687988 pi
 12'b010110000010: begin out_real=16'b1101110001001000; out_imag=16'b0011010100011011; end // in_theta = 0.688477 pi
 12'b010110000011: begin out_real=16'b1101110000110011; out_imag=16'b0011010100001101; end // in_theta = 0.688965 pi
 12'b010110000100: begin out_real=16'b1101110000011110; out_imag=16'b0011010011111111; end // in_theta = 0.689453 pi
 12'b010110000101: begin out_real=16'b1101110000001001; out_imag=16'b0011010011110001; end // in_theta = 0.689941 pi
 12'b010110000110: begin out_real=16'b1101101111110101; out_imag=16'b0011010011100010; end // in_theta = 0.690430 pi
 12'b010110000111: begin out_real=16'b1101101111100000; out_imag=16'b0011010011010100; end // in_theta = 0.690918 pi
 12'b010110001000: begin out_real=16'b1101101111001011; out_imag=16'b0011010011000110; end // in_theta = 0.691406 pi
 12'b010110001001: begin out_real=16'b1101101110110110; out_imag=16'b0011010010111000; end // in_theta = 0.691895 pi
 12'b010110001010: begin out_real=16'b1101101110100010; out_imag=16'b0011010010101010; end // in_theta = 0.692383 pi
 12'b010110001011: begin out_real=16'b1101101110001101; out_imag=16'b0011010010011011; end // in_theta = 0.692871 pi
 12'b010110001100: begin out_real=16'b1101101101111000; out_imag=16'b0011010010001101; end // in_theta = 0.693359 pi
 12'b010110001101: begin out_real=16'b1101101101100100; out_imag=16'b0011010001111111; end // in_theta = 0.693848 pi
 12'b010110001110: begin out_real=16'b1101101101001111; out_imag=16'b0011010001110000; end // in_theta = 0.694336 pi
 12'b010110001111: begin out_real=16'b1101101100111011; out_imag=16'b0011010001100010; end // in_theta = 0.694824 pi
 12'b010110010000: begin out_real=16'b1101101100100110; out_imag=16'b0011010001010011; end // in_theta = 0.695313 pi
 12'b010110010001: begin out_real=16'b1101101100010001; out_imag=16'b0011010001000101; end // in_theta = 0.695801 pi
 12'b010110010010: begin out_real=16'b1101101011111101; out_imag=16'b0011010000110110; end // in_theta = 0.696289 pi
 12'b010110010011: begin out_real=16'b1101101011101000; out_imag=16'b0011010000101000; end // in_theta = 0.696777 pi
 12'b010110010100: begin out_real=16'b1101101011010100; out_imag=16'b0011010000011001; end // in_theta = 0.697266 pi
 12'b010110010101: begin out_real=16'b1101101010111111; out_imag=16'b0011010000001011; end // in_theta = 0.697754 pi
 12'b010110010110: begin out_real=16'b1101101010101011; out_imag=16'b0011001111111100; end // in_theta = 0.698242 pi
 12'b010110010111: begin out_real=16'b1101101010010111; out_imag=16'b0011001111101101; end // in_theta = 0.698730 pi
 12'b010110011000: begin out_real=16'b1101101010000010; out_imag=16'b0011001111011111; end // in_theta = 0.699219 pi
 12'b010110011001: begin out_real=16'b1101101001101110; out_imag=16'b0011001111010000; end // in_theta = 0.699707 pi
 12'b010110011010: begin out_real=16'b1101101001011010; out_imag=16'b0011001111000001; end // in_theta = 0.700195 pi
 12'b010110011011: begin out_real=16'b1101101001000101; out_imag=16'b0011001110110010; end // in_theta = 0.700684 pi
 12'b010110011100: begin out_real=16'b1101101000110001; out_imag=16'b0011001110100011; end // in_theta = 0.701172 pi
 12'b010110011101: begin out_real=16'b1101101000011101; out_imag=16'b0011001110010101; end // in_theta = 0.701660 pi
 12'b010110011110: begin out_real=16'b1101101000001000; out_imag=16'b0011001110000110; end // in_theta = 0.702148 pi
 12'b010110011111: begin out_real=16'b1101100111110100; out_imag=16'b0011001101110111; end // in_theta = 0.702637 pi
 12'b010110100000: begin out_real=16'b1101100111100000; out_imag=16'b0011001101101000; end // in_theta = 0.703125 pi
 12'b010110100001: begin out_real=16'b1101100111001100; out_imag=16'b0011001101011001; end // in_theta = 0.703613 pi
 12'b010110100010: begin out_real=16'b1101100110111000; out_imag=16'b0011001101001010; end // in_theta = 0.704102 pi
 12'b010110100011: begin out_real=16'b1101100110100100; out_imag=16'b0011001100111011; end // in_theta = 0.704590 pi
 12'b010110100100: begin out_real=16'b1101100110001111; out_imag=16'b0011001100101100; end // in_theta = 0.705078 pi
 12'b010110100101: begin out_real=16'b1101100101111011; out_imag=16'b0011001100011101; end // in_theta = 0.705566 pi
 12'b010110100110: begin out_real=16'b1101100101100111; out_imag=16'b0011001100001101; end // in_theta = 0.706055 pi
 12'b010110100111: begin out_real=16'b1101100101010011; out_imag=16'b0011001011111110; end // in_theta = 0.706543 pi
 12'b010110101000: begin out_real=16'b1101100100111111; out_imag=16'b0011001011101111; end // in_theta = 0.707031 pi
 12'b010110101001: begin out_real=16'b1101100100101011; out_imag=16'b0011001011100000; end // in_theta = 0.707520 pi
 12'b010110101010: begin out_real=16'b1101100100010111; out_imag=16'b0011001011010000; end // in_theta = 0.708008 pi
 12'b010110101011: begin out_real=16'b1101100100000011; out_imag=16'b0011001011000001; end // in_theta = 0.708496 pi
 12'b010110101100: begin out_real=16'b1101100011101111; out_imag=16'b0011001010110010; end // in_theta = 0.708984 pi
 12'b010110101101: begin out_real=16'b1101100011011100; out_imag=16'b0011001010100011; end // in_theta = 0.709473 pi
 12'b010110101110: begin out_real=16'b1101100011001000; out_imag=16'b0011001010010011; end // in_theta = 0.709961 pi
 12'b010110101111: begin out_real=16'b1101100010110100; out_imag=16'b0011001010000100; end // in_theta = 0.710449 pi
 12'b010110110000: begin out_real=16'b1101100010100000; out_imag=16'b0011001001110100; end // in_theta = 0.710938 pi
 12'b010110110001: begin out_real=16'b1101100010001100; out_imag=16'b0011001001100101; end // in_theta = 0.711426 pi
 12'b010110110010: begin out_real=16'b1101100001111000; out_imag=16'b0011001001010101; end // in_theta = 0.711914 pi
 12'b010110110011: begin out_real=16'b1101100001100101; out_imag=16'b0011001001000110; end // in_theta = 0.712402 pi
 12'b010110110100: begin out_real=16'b1101100001010001; out_imag=16'b0011001000110110; end // in_theta = 0.712891 pi
 12'b010110110101: begin out_real=16'b1101100000111101; out_imag=16'b0011001000100111; end // in_theta = 0.713379 pi
 12'b010110110110: begin out_real=16'b1101100000101010; out_imag=16'b0011001000010111; end // in_theta = 0.713867 pi
 12'b010110110111: begin out_real=16'b1101100000010110; out_imag=16'b0011001000000111; end // in_theta = 0.714355 pi
 12'b010110111000: begin out_real=16'b1101100000000010; out_imag=16'b0011000111111000; end // in_theta = 0.714844 pi
 12'b010110111001: begin out_real=16'b1101011111101111; out_imag=16'b0011000111101000; end // in_theta = 0.715332 pi
 12'b010110111010: begin out_real=16'b1101011111011011; out_imag=16'b0011000111011000; end // in_theta = 0.715820 pi
 12'b010110111011: begin out_real=16'b1101011111001000; out_imag=16'b0011000111001000; end // in_theta = 0.716309 pi
 12'b010110111100: begin out_real=16'b1101011110110100; out_imag=16'b0011000110111001; end // in_theta = 0.716797 pi
 12'b010110111101: begin out_real=16'b1101011110100000; out_imag=16'b0011000110101001; end // in_theta = 0.717285 pi
 12'b010110111110: begin out_real=16'b1101011110001101; out_imag=16'b0011000110011001; end // in_theta = 0.717773 pi
 12'b010110111111: begin out_real=16'b1101011101111010; out_imag=16'b0011000110001001; end // in_theta = 0.718262 pi
 12'b010111000000: begin out_real=16'b1101011101100110; out_imag=16'b0011000101111001; end // in_theta = 0.718750 pi
 12'b010111000001: begin out_real=16'b1101011101010011; out_imag=16'b0011000101101001; end // in_theta = 0.719238 pi
 12'b010111000010: begin out_real=16'b1101011100111111; out_imag=16'b0011000101011001; end // in_theta = 0.719727 pi
 12'b010111000011: begin out_real=16'b1101011100101100; out_imag=16'b0011000101001001; end // in_theta = 0.720215 pi
 12'b010111000100: begin out_real=16'b1101011100011001; out_imag=16'b0011000100111001; end // in_theta = 0.720703 pi
 12'b010111000101: begin out_real=16'b1101011100000101; out_imag=16'b0011000100101001; end // in_theta = 0.721191 pi
 12'b010111000110: begin out_real=16'b1101011011110010; out_imag=16'b0011000100011001; end // in_theta = 0.721680 pi
 12'b010111000111: begin out_real=16'b1101011011011111; out_imag=16'b0011000100001001; end // in_theta = 0.722168 pi
 12'b010111001000: begin out_real=16'b1101011011001011; out_imag=16'b0011000011111001; end // in_theta = 0.722656 pi
 12'b010111001001: begin out_real=16'b1101011010111000; out_imag=16'b0011000011101000; end // in_theta = 0.723145 pi
 12'b010111001010: begin out_real=16'b1101011010100101; out_imag=16'b0011000011011000; end // in_theta = 0.723633 pi
 12'b010111001011: begin out_real=16'b1101011010010010; out_imag=16'b0011000011001000; end // in_theta = 0.724121 pi
 12'b010111001100: begin out_real=16'b1101011001111111; out_imag=16'b0011000010111000; end // in_theta = 0.724609 pi
 12'b010111001101: begin out_real=16'b1101011001101100; out_imag=16'b0011000010100111; end // in_theta = 0.725098 pi
 12'b010111001110: begin out_real=16'b1101011001011001; out_imag=16'b0011000010010111; end // in_theta = 0.725586 pi
 12'b010111001111: begin out_real=16'b1101011001000101; out_imag=16'b0011000010000111; end // in_theta = 0.726074 pi
 12'b010111010000: begin out_real=16'b1101011000110010; out_imag=16'b0011000001110110; end // in_theta = 0.726562 pi
 12'b010111010001: begin out_real=16'b1101011000011111; out_imag=16'b0011000001100110; end // in_theta = 0.727051 pi
 12'b010111010010: begin out_real=16'b1101011000001100; out_imag=16'b0011000001010101; end // in_theta = 0.727539 pi
 12'b010111010011: begin out_real=16'b1101010111111001; out_imag=16'b0011000001000101; end // in_theta = 0.728027 pi
 12'b010111010100: begin out_real=16'b1101010111100110; out_imag=16'b0011000000110100; end // in_theta = 0.728516 pi
 12'b010111010101: begin out_real=16'b1101010111010100; out_imag=16'b0011000000100100; end // in_theta = 0.729004 pi
 12'b010111010110: begin out_real=16'b1101010111000001; out_imag=16'b0011000000010011; end // in_theta = 0.729492 pi
 12'b010111010111: begin out_real=16'b1101010110101110; out_imag=16'b0011000000000010; end // in_theta = 0.729980 pi
 12'b010111011000: begin out_real=16'b1101010110011011; out_imag=16'b0010111111110010; end // in_theta = 0.730469 pi
 12'b010111011001: begin out_real=16'b1101010110001000; out_imag=16'b0010111111100001; end // in_theta = 0.730957 pi
 12'b010111011010: begin out_real=16'b1101010101110101; out_imag=16'b0010111111010000; end // in_theta = 0.731445 pi
 12'b010111011011: begin out_real=16'b1101010101100011; out_imag=16'b0010111111000000; end // in_theta = 0.731934 pi
 12'b010111011100: begin out_real=16'b1101010101010000; out_imag=16'b0010111110101111; end // in_theta = 0.732422 pi
 12'b010111011101: begin out_real=16'b1101010100111101; out_imag=16'b0010111110011110; end // in_theta = 0.732910 pi
 12'b010111011110: begin out_real=16'b1101010100101010; out_imag=16'b0010111110001101; end // in_theta = 0.733398 pi
 12'b010111011111: begin out_real=16'b1101010100011000; out_imag=16'b0010111101111101; end // in_theta = 0.733887 pi
 12'b010111100000: begin out_real=16'b1101010100000101; out_imag=16'b0010111101101100; end // in_theta = 0.734375 pi
 12'b010111100001: begin out_real=16'b1101010011110011; out_imag=16'b0010111101011011; end // in_theta = 0.734863 pi
 12'b010111100010: begin out_real=16'b1101010011100000; out_imag=16'b0010111101001010; end // in_theta = 0.735352 pi
 12'b010111100011: begin out_real=16'b1101010011001101; out_imag=16'b0010111100111001; end // in_theta = 0.735840 pi
 12'b010111100100: begin out_real=16'b1101010010111011; out_imag=16'b0010111100101000; end // in_theta = 0.736328 pi
 12'b010111100101: begin out_real=16'b1101010010101000; out_imag=16'b0010111100010111; end // in_theta = 0.736816 pi
 12'b010111100110: begin out_real=16'b1101010010010110; out_imag=16'b0010111100000110; end // in_theta = 0.737305 pi
 12'b010111100111: begin out_real=16'b1101010010000011; out_imag=16'b0010111011110101; end // in_theta = 0.737793 pi
 12'b010111101000: begin out_real=16'b1101010001110001; out_imag=16'b0010111011100100; end // in_theta = 0.738281 pi
 12'b010111101001: begin out_real=16'b1101010001011111; out_imag=16'b0010111011010011; end // in_theta = 0.738770 pi
 12'b010111101010: begin out_real=16'b1101010001001100; out_imag=16'b0010111011000010; end // in_theta = 0.739258 pi
 12'b010111101011: begin out_real=16'b1101010000111010; out_imag=16'b0010111010110000; end // in_theta = 0.739746 pi
 12'b010111101100: begin out_real=16'b1101010000101000; out_imag=16'b0010111010011111; end // in_theta = 0.740234 pi
 12'b010111101101: begin out_real=16'b1101010000010101; out_imag=16'b0010111010001110; end // in_theta = 0.740723 pi
 12'b010111101110: begin out_real=16'b1101010000000011; out_imag=16'b0010111001111101; end // in_theta = 0.741211 pi
 12'b010111101111: begin out_real=16'b1101001111110001; out_imag=16'b0010111001101011; end // in_theta = 0.741699 pi
 12'b010111110000: begin out_real=16'b1101001111011111; out_imag=16'b0010111001011010; end // in_theta = 0.742188 pi
 12'b010111110001: begin out_real=16'b1101001111001100; out_imag=16'b0010111001001001; end // in_theta = 0.742676 pi
 12'b010111110010: begin out_real=16'b1101001110111010; out_imag=16'b0010111000110111; end // in_theta = 0.743164 pi
 12'b010111110011: begin out_real=16'b1101001110101000; out_imag=16'b0010111000100110; end // in_theta = 0.743652 pi
 12'b010111110100: begin out_real=16'b1101001110010110; out_imag=16'b0010111000010101; end // in_theta = 0.744141 pi
 12'b010111110101: begin out_real=16'b1101001110000100; out_imag=16'b0010111000000011; end // in_theta = 0.744629 pi
 12'b010111110110: begin out_real=16'b1101001101110010; out_imag=16'b0010110111110010; end // in_theta = 0.745117 pi
 12'b010111110111: begin out_real=16'b1101001101100000; out_imag=16'b0010110111100000; end // in_theta = 0.745605 pi
 12'b010111111000: begin out_real=16'b1101001101001110; out_imag=16'b0010110111001111; end // in_theta = 0.746094 pi
 12'b010111111001: begin out_real=16'b1101001100111100; out_imag=16'b0010110110111101; end // in_theta = 0.746582 pi
 12'b010111111010: begin out_real=16'b1101001100101010; out_imag=16'b0010110110101011; end // in_theta = 0.747070 pi
 12'b010111111011: begin out_real=16'b1101001100011000; out_imag=16'b0010110110011010; end // in_theta = 0.747559 pi
 12'b010111111100: begin out_real=16'b1101001100000110; out_imag=16'b0010110110001000; end // in_theta = 0.748047 pi
 12'b010111111101: begin out_real=16'b1101001011110100; out_imag=16'b0010110101110110; end // in_theta = 0.748535 pi
 12'b010111111110: begin out_real=16'b1101001011100010; out_imag=16'b0010110101100101; end // in_theta = 0.749023 pi
 12'b010111111111: begin out_real=16'b1101001011010001; out_imag=16'b0010110101010011; end // in_theta = 0.749512 pi
 12'b011000000000: begin out_real=16'b1101001010111111; out_imag=16'b0010110101000001; end // in_theta = 0.750000 pi
 12'b011000000001: begin out_real=16'b1101001010101101; out_imag=16'b0010110100101111; end // in_theta = 0.750488 pi
 12'b011000000010: begin out_real=16'b1101001010011011; out_imag=16'b0010110100011110; end // in_theta = 0.750977 pi
 12'b011000000011: begin out_real=16'b1101001010001010; out_imag=16'b0010110100001100; end // in_theta = 0.751465 pi
 12'b011000000100: begin out_real=16'b1101001001111000; out_imag=16'b0010110011111010; end // in_theta = 0.751953 pi
 12'b011000000101: begin out_real=16'b1101001001100110; out_imag=16'b0010110011101000; end // in_theta = 0.752441 pi
 12'b011000000110: begin out_real=16'b1101001001010101; out_imag=16'b0010110011010110; end // in_theta = 0.752930 pi
 12'b011000000111: begin out_real=16'b1101001001000011; out_imag=16'b0010110011000100; end // in_theta = 0.753418 pi
 12'b011000001000: begin out_real=16'b1101001000110001; out_imag=16'b0010110010110010; end // in_theta = 0.753906 pi
 12'b011000001001: begin out_real=16'b1101001000100000; out_imag=16'b0010110010100000; end // in_theta = 0.754395 pi
 12'b011000001010: begin out_real=16'b1101001000001110; out_imag=16'b0010110010001110; end // in_theta = 0.754883 pi
 12'b011000001011: begin out_real=16'b1101000111111101; out_imag=16'b0010110001111100; end // in_theta = 0.755371 pi
 12'b011000001100: begin out_real=16'b1101000111101011; out_imag=16'b0010110001101010; end // in_theta = 0.755859 pi
 12'b011000001101: begin out_real=16'b1101000111011010; out_imag=16'b0010110001011000; end // in_theta = 0.756348 pi
 12'b011000001110: begin out_real=16'b1101000111001001; out_imag=16'b0010110001000110; end // in_theta = 0.756836 pi
 12'b011000001111: begin out_real=16'b1101000110110111; out_imag=16'b0010110000110100; end // in_theta = 0.757324 pi
 12'b011000010000: begin out_real=16'b1101000110100110; out_imag=16'b0010110000100001; end // in_theta = 0.757813 pi
 12'b011000010001: begin out_real=16'b1101000110010101; out_imag=16'b0010110000001111; end // in_theta = 0.758301 pi
 12'b011000010010: begin out_real=16'b1101000110000011; out_imag=16'b0010101111111101; end // in_theta = 0.758789 pi
 12'b011000010011: begin out_real=16'b1101000101110010; out_imag=16'b0010101111101011; end // in_theta = 0.759277 pi
 12'b011000010100: begin out_real=16'b1101000101100001; out_imag=16'b0010101111011000; end // in_theta = 0.759766 pi
 12'b011000010101: begin out_real=16'b1101000101010000; out_imag=16'b0010101111000110; end // in_theta = 0.760254 pi
 12'b011000010110: begin out_real=16'b1101000100111110; out_imag=16'b0010101110110100; end // in_theta = 0.760742 pi
 12'b011000010111: begin out_real=16'b1101000100101101; out_imag=16'b0010101110100001; end // in_theta = 0.761230 pi
 12'b011000011000: begin out_real=16'b1101000100011100; out_imag=16'b0010101110001111; end // in_theta = 0.761719 pi
 12'b011000011001: begin out_real=16'b1101000100001011; out_imag=16'b0010101101111101; end // in_theta = 0.762207 pi
 12'b011000011010: begin out_real=16'b1101000011111010; out_imag=16'b0010101101101010; end // in_theta = 0.762695 pi
 12'b011000011011: begin out_real=16'b1101000011101001; out_imag=16'b0010101101011000; end // in_theta = 0.763184 pi
 12'b011000011100: begin out_real=16'b1101000011011000; out_imag=16'b0010101101000101; end // in_theta = 0.763672 pi
 12'b011000011101: begin out_real=16'b1101000011000111; out_imag=16'b0010101100110011; end // in_theta = 0.764160 pi
 12'b011000011110: begin out_real=16'b1101000010110110; out_imag=16'b0010101100100000; end // in_theta = 0.764648 pi
 12'b011000011111: begin out_real=16'b1101000010100101; out_imag=16'b0010101100001101; end // in_theta = 0.765137 pi
 12'b011000100000: begin out_real=16'b1101000010010100; out_imag=16'b0010101011111011; end // in_theta = 0.765625 pi
 12'b011000100001: begin out_real=16'b1101000010000011; out_imag=16'b0010101011101000; end // in_theta = 0.766113 pi
 12'b011000100010: begin out_real=16'b1101000001110011; out_imag=16'b0010101011010110; end // in_theta = 0.766602 pi
 12'b011000100011: begin out_real=16'b1101000001100010; out_imag=16'b0010101011000011; end // in_theta = 0.767090 pi
 12'b011000100100: begin out_real=16'b1101000001010001; out_imag=16'b0010101010110000; end // in_theta = 0.767578 pi
 12'b011000100101: begin out_real=16'b1101000001000000; out_imag=16'b0010101010011101; end // in_theta = 0.768066 pi
 12'b011000100110: begin out_real=16'b1101000000110000; out_imag=16'b0010101010001011; end // in_theta = 0.768555 pi
 12'b011000100111: begin out_real=16'b1101000000011111; out_imag=16'b0010101001111000; end // in_theta = 0.769043 pi
 12'b011000101000: begin out_real=16'b1101000000001110; out_imag=16'b0010101001100101; end // in_theta = 0.769531 pi
 12'b011000101001: begin out_real=16'b1100111111111110; out_imag=16'b0010101001010010; end // in_theta = 0.770020 pi
 12'b011000101010: begin out_real=16'b1100111111101101; out_imag=16'b0010101000111111; end // in_theta = 0.770508 pi
 12'b011000101011: begin out_real=16'b1100111111011100; out_imag=16'b0010101000101100; end // in_theta = 0.770996 pi
 12'b011000101100: begin out_real=16'b1100111111001100; out_imag=16'b0010101000011010; end // in_theta = 0.771484 pi
 12'b011000101101: begin out_real=16'b1100111110111011; out_imag=16'b0010101000000111; end // in_theta = 0.771973 pi
 12'b011000101110: begin out_real=16'b1100111110101011; out_imag=16'b0010100111110100; end // in_theta = 0.772461 pi
 12'b011000101111: begin out_real=16'b1100111110011010; out_imag=16'b0010100111100001; end // in_theta = 0.772949 pi
 12'b011000110000: begin out_real=16'b1100111110001010; out_imag=16'b0010100111001110; end // in_theta = 0.773438 pi
 12'b011000110001: begin out_real=16'b1100111101111001; out_imag=16'b0010100110111011; end // in_theta = 0.773926 pi
 12'b011000110010: begin out_real=16'b1100111101101001; out_imag=16'b0010100110100111; end // in_theta = 0.774414 pi
 12'b011000110011: begin out_real=16'b1100111101011001; out_imag=16'b0010100110010100; end // in_theta = 0.774902 pi
 12'b011000110100: begin out_real=16'b1100111101001000; out_imag=16'b0010100110000001; end // in_theta = 0.775391 pi
 12'b011000110101: begin out_real=16'b1100111100111000; out_imag=16'b0010100101101110; end // in_theta = 0.775879 pi
 12'b011000110110: begin out_real=16'b1100111100101000; out_imag=16'b0010100101011011; end // in_theta = 0.776367 pi
 12'b011000110111: begin out_real=16'b1100111100011000; out_imag=16'b0010100101001000; end // in_theta = 0.776855 pi
 12'b011000111000: begin out_real=16'b1100111100000111; out_imag=16'b0010100100110101; end // in_theta = 0.777344 pi
 12'b011000111001: begin out_real=16'b1100111011110111; out_imag=16'b0010100100100001; end // in_theta = 0.777832 pi
 12'b011000111010: begin out_real=16'b1100111011100111; out_imag=16'b0010100100001110; end // in_theta = 0.778320 pi
 12'b011000111011: begin out_real=16'b1100111011010111; out_imag=16'b0010100011111011; end // in_theta = 0.778809 pi
 12'b011000111100: begin out_real=16'b1100111011000111; out_imag=16'b0010100011100111; end // in_theta = 0.779297 pi
 12'b011000111101: begin out_real=16'b1100111010110111; out_imag=16'b0010100011010100; end // in_theta = 0.779785 pi
 12'b011000111110: begin out_real=16'b1100111010100111; out_imag=16'b0010100011000001; end // in_theta = 0.780273 pi
 12'b011000111111: begin out_real=16'b1100111010010111; out_imag=16'b0010100010101101; end // in_theta = 0.780762 pi
 12'b011001000000: begin out_real=16'b1100111010000111; out_imag=16'b0010100010011010; end // in_theta = 0.781250 pi
 12'b011001000001: begin out_real=16'b1100111001110111; out_imag=16'b0010100010000110; end // in_theta = 0.781738 pi
 12'b011001000010: begin out_real=16'b1100111001100111; out_imag=16'b0010100001110011; end // in_theta = 0.782227 pi
 12'b011001000011: begin out_real=16'b1100111001010111; out_imag=16'b0010100001100000; end // in_theta = 0.782715 pi
 12'b011001000100: begin out_real=16'b1100111001000111; out_imag=16'b0010100001001100; end // in_theta = 0.783203 pi
 12'b011001000101: begin out_real=16'b1100111000111000; out_imag=16'b0010100000111000; end // in_theta = 0.783691 pi
 12'b011001000110: begin out_real=16'b1100111000101000; out_imag=16'b0010100000100101; end // in_theta = 0.784180 pi
 12'b011001000111: begin out_real=16'b1100111000011000; out_imag=16'b0010100000010001; end // in_theta = 0.784668 pi
 12'b011001001000: begin out_real=16'b1100111000001000; out_imag=16'b0010011111111110; end // in_theta = 0.785156 pi
 12'b011001001001: begin out_real=16'b1100110111111001; out_imag=16'b0010011111101010; end // in_theta = 0.785645 pi
 12'b011001001010: begin out_real=16'b1100110111101001; out_imag=16'b0010011111010110; end // in_theta = 0.786133 pi
 12'b011001001011: begin out_real=16'b1100110111011001; out_imag=16'b0010011111000011; end // in_theta = 0.786621 pi
 12'b011001001100: begin out_real=16'b1100110111001010; out_imag=16'b0010011110101111; end // in_theta = 0.787109 pi
 12'b011001001101: begin out_real=16'b1100110110111010; out_imag=16'b0010011110011011; end // in_theta = 0.787598 pi
 12'b011001001110: begin out_real=16'b1100110110101011; out_imag=16'b0010011110001000; end // in_theta = 0.788086 pi
 12'b011001001111: begin out_real=16'b1100110110011011; out_imag=16'b0010011101110100; end // in_theta = 0.788574 pi
 12'b011001010000: begin out_real=16'b1100110110001100; out_imag=16'b0010011101100000; end // in_theta = 0.789063 pi
 12'b011001010001: begin out_real=16'b1100110101111100; out_imag=16'b0010011101001100; end // in_theta = 0.789551 pi
 12'b011001010010: begin out_real=16'b1100110101101101; out_imag=16'b0010011100111000; end // in_theta = 0.790039 pi
 12'b011001010011: begin out_real=16'b1100110101011101; out_imag=16'b0010011100100100; end // in_theta = 0.790527 pi
 12'b011001010100: begin out_real=16'b1100110101001110; out_imag=16'b0010011100010001; end // in_theta = 0.791016 pi
 12'b011001010101: begin out_real=16'b1100110100111111; out_imag=16'b0010011011111101; end // in_theta = 0.791504 pi
 12'b011001010110: begin out_real=16'b1100110100110000; out_imag=16'b0010011011101001; end // in_theta = 0.791992 pi
 12'b011001010111: begin out_real=16'b1100110100100000; out_imag=16'b0010011011010101; end // in_theta = 0.792480 pi
 12'b011001011000: begin out_real=16'b1100110100010001; out_imag=16'b0010011011000001; end // in_theta = 0.792969 pi
 12'b011001011001: begin out_real=16'b1100110100000010; out_imag=16'b0010011010101101; end // in_theta = 0.793457 pi
 12'b011001011010: begin out_real=16'b1100110011110011; out_imag=16'b0010011010011001; end // in_theta = 0.793945 pi
 12'b011001011011: begin out_real=16'b1100110011100011; out_imag=16'b0010011010000101; end // in_theta = 0.794434 pi
 12'b011001011100: begin out_real=16'b1100110011010100; out_imag=16'b0010011001110001; end // in_theta = 0.794922 pi
 12'b011001011101: begin out_real=16'b1100110011000101; out_imag=16'b0010011001011100; end // in_theta = 0.795410 pi
 12'b011001011110: begin out_real=16'b1100110010110110; out_imag=16'b0010011001001000; end // in_theta = 0.795898 pi
 12'b011001011111: begin out_real=16'b1100110010100111; out_imag=16'b0010011000110100; end // in_theta = 0.796387 pi
 12'b011001100000: begin out_real=16'b1100110010011000; out_imag=16'b0010011000100000; end // in_theta = 0.796875 pi
 12'b011001100001: begin out_real=16'b1100110010001001; out_imag=16'b0010011000001100; end // in_theta = 0.797363 pi
 12'b011001100010: begin out_real=16'b1100110001111010; out_imag=16'b0010010111111000; end // in_theta = 0.797852 pi
 12'b011001100011: begin out_real=16'b1100110001101011; out_imag=16'b0010010111100011; end // in_theta = 0.798340 pi
 12'b011001100100: begin out_real=16'b1100110001011101; out_imag=16'b0010010111001111; end // in_theta = 0.798828 pi
 12'b011001100101: begin out_real=16'b1100110001001110; out_imag=16'b0010010110111011; end // in_theta = 0.799316 pi
 12'b011001100110: begin out_real=16'b1100110000111111; out_imag=16'b0010010110100110; end // in_theta = 0.799805 pi
 12'b011001100111: begin out_real=16'b1100110000110000; out_imag=16'b0010010110010010; end // in_theta = 0.800293 pi
 12'b011001101000: begin out_real=16'b1100110000100001; out_imag=16'b0010010101111110; end // in_theta = 0.800781 pi
 12'b011001101001: begin out_real=16'b1100110000010011; out_imag=16'b0010010101101001; end // in_theta = 0.801270 pi
 12'b011001101010: begin out_real=16'b1100110000000100; out_imag=16'b0010010101010101; end // in_theta = 0.801758 pi
 12'b011001101011: begin out_real=16'b1100101111110101; out_imag=16'b0010010101000001; end // in_theta = 0.802246 pi
 12'b011001101100: begin out_real=16'b1100101111100111; out_imag=16'b0010010100101100; end // in_theta = 0.802734 pi
 12'b011001101101: begin out_real=16'b1100101111011000; out_imag=16'b0010010100011000; end // in_theta = 0.803223 pi
 12'b011001101110: begin out_real=16'b1100101111001010; out_imag=16'b0010010100000011; end // in_theta = 0.803711 pi
 12'b011001101111: begin out_real=16'b1100101110111011; out_imag=16'b0010010011101111; end // in_theta = 0.804199 pi
 12'b011001110000: begin out_real=16'b1100101110101101; out_imag=16'b0010010011011010; end // in_theta = 0.804688 pi
 12'b011001110001: begin out_real=16'b1100101110011110; out_imag=16'b0010010011000101; end // in_theta = 0.805176 pi
 12'b011001110010: begin out_real=16'b1100101110010000; out_imag=16'b0010010010110001; end // in_theta = 0.805664 pi
 12'b011001110011: begin out_real=16'b1100101110000001; out_imag=16'b0010010010011100; end // in_theta = 0.806152 pi
 12'b011001110100: begin out_real=16'b1100101101110011; out_imag=16'b0010010010001000; end // in_theta = 0.806641 pi
 12'b011001110101: begin out_real=16'b1100101101100101; out_imag=16'b0010010001110011; end // in_theta = 0.807129 pi
 12'b011001110110: begin out_real=16'b1100101101010110; out_imag=16'b0010010001011110; end // in_theta = 0.807617 pi
 12'b011001110111: begin out_real=16'b1100101101001000; out_imag=16'b0010010001001010; end // in_theta = 0.808105 pi
 12'b011001111000: begin out_real=16'b1100101100111010; out_imag=16'b0010010000110101; end // in_theta = 0.808594 pi
 12'b011001111001: begin out_real=16'b1100101100101100; out_imag=16'b0010010000100000; end // in_theta = 0.809082 pi
 12'b011001111010: begin out_real=16'b1100101100011110; out_imag=16'b0010010000001011; end // in_theta = 0.809570 pi
 12'b011001111011: begin out_real=16'b1100101100001111; out_imag=16'b0010001111110111; end // in_theta = 0.810059 pi
 12'b011001111100: begin out_real=16'b1100101100000001; out_imag=16'b0010001111100010; end // in_theta = 0.810547 pi
 12'b011001111101: begin out_real=16'b1100101011110011; out_imag=16'b0010001111001101; end // in_theta = 0.811035 pi
 12'b011001111110: begin out_real=16'b1100101011100101; out_imag=16'b0010001110111000; end // in_theta = 0.811523 pi
 12'b011001111111: begin out_real=16'b1100101011010111; out_imag=16'b0010001110100011; end // in_theta = 0.812012 pi
 12'b011010000000: begin out_real=16'b1100101011001001; out_imag=16'b0010001110001110; end // in_theta = 0.812500 pi
 12'b011010000001: begin out_real=16'b1100101010111011; out_imag=16'b0010001101111010; end // in_theta = 0.812988 pi
 12'b011010000010: begin out_real=16'b1100101010101101; out_imag=16'b0010001101100101; end // in_theta = 0.813477 pi
 12'b011010000011: begin out_real=16'b1100101010011111; out_imag=16'b0010001101010000; end // in_theta = 0.813965 pi
 12'b011010000100: begin out_real=16'b1100101010010010; out_imag=16'b0010001100111011; end // in_theta = 0.814453 pi
 12'b011010000101: begin out_real=16'b1100101010000100; out_imag=16'b0010001100100110; end // in_theta = 0.814941 pi
 12'b011010000110: begin out_real=16'b1100101001110110; out_imag=16'b0010001100010001; end // in_theta = 0.815430 pi
 12'b011010000111: begin out_real=16'b1100101001101000; out_imag=16'b0010001011111100; end // in_theta = 0.815918 pi
 12'b011010001000: begin out_real=16'b1100101001011011; out_imag=16'b0010001011100111; end // in_theta = 0.816406 pi
 12'b011010001001: begin out_real=16'b1100101001001101; out_imag=16'b0010001011010010; end // in_theta = 0.816895 pi
 12'b011010001010: begin out_real=16'b1100101000111111; out_imag=16'b0010001010111100; end // in_theta = 0.817383 pi
 12'b011010001011: begin out_real=16'b1100101000110010; out_imag=16'b0010001010100111; end // in_theta = 0.817871 pi
 12'b011010001100: begin out_real=16'b1100101000100100; out_imag=16'b0010001010010010; end // in_theta = 0.818359 pi
 12'b011010001101: begin out_real=16'b1100101000010110; out_imag=16'b0010001001111101; end // in_theta = 0.818848 pi
 12'b011010001110: begin out_real=16'b1100101000001001; out_imag=16'b0010001001101000; end // in_theta = 0.819336 pi
 12'b011010001111: begin out_real=16'b1100100111111011; out_imag=16'b0010001001010011; end // in_theta = 0.819824 pi
 12'b011010010000: begin out_real=16'b1100100111101110; out_imag=16'b0010001000111101; end // in_theta = 0.820313 pi
 12'b011010010001: begin out_real=16'b1100100111100000; out_imag=16'b0010001000101000; end // in_theta = 0.820801 pi
 12'b011010010010: begin out_real=16'b1100100111010011; out_imag=16'b0010001000010011; end // in_theta = 0.821289 pi
 12'b011010010011: begin out_real=16'b1100100111000110; out_imag=16'b0010000111111110; end // in_theta = 0.821777 pi
 12'b011010010100: begin out_real=16'b1100100110111000; out_imag=16'b0010000111101000; end // in_theta = 0.822266 pi
 12'b011010010101: begin out_real=16'b1100100110101011; out_imag=16'b0010000111010011; end // in_theta = 0.822754 pi
 12'b011010010110: begin out_real=16'b1100100110011110; out_imag=16'b0010000110111110; end // in_theta = 0.823242 pi
 12'b011010010111: begin out_real=16'b1100100110010001; out_imag=16'b0010000110101000; end // in_theta = 0.823730 pi
 12'b011010011000: begin out_real=16'b1100100110000011; out_imag=16'b0010000110010011; end // in_theta = 0.824219 pi
 12'b011010011001: begin out_real=16'b1100100101110110; out_imag=16'b0010000101111101; end // in_theta = 0.824707 pi
 12'b011010011010: begin out_real=16'b1100100101101001; out_imag=16'b0010000101101000; end // in_theta = 0.825195 pi
 12'b011010011011: begin out_real=16'b1100100101011100; out_imag=16'b0010000101010011; end // in_theta = 0.825684 pi
 12'b011010011100: begin out_real=16'b1100100101001111; out_imag=16'b0010000100111101; end // in_theta = 0.826172 pi
 12'b011010011101: begin out_real=16'b1100100101000010; out_imag=16'b0010000100101000; end // in_theta = 0.826660 pi
 12'b011010011110: begin out_real=16'b1100100100110101; out_imag=16'b0010000100010010; end // in_theta = 0.827148 pi
 12'b011010011111: begin out_real=16'b1100100100101000; out_imag=16'b0010000011111101; end // in_theta = 0.827637 pi
 12'b011010100000: begin out_real=16'b1100100100011011; out_imag=16'b0010000011100111; end // in_theta = 0.828125 pi
 12'b011010100001: begin out_real=16'b1100100100001110; out_imag=16'b0010000011010001; end // in_theta = 0.828613 pi
 12'b011010100010: begin out_real=16'b1100100100000001; out_imag=16'b0010000010111100; end // in_theta = 0.829102 pi
 12'b011010100011: begin out_real=16'b1100100011110100; out_imag=16'b0010000010100110; end // in_theta = 0.829590 pi
 12'b011010100100: begin out_real=16'b1100100011101000; out_imag=16'b0010000010010001; end // in_theta = 0.830078 pi
 12'b011010100101: begin out_real=16'b1100100011011011; out_imag=16'b0010000001111011; end // in_theta = 0.830566 pi
 12'b011010100110: begin out_real=16'b1100100011001110; out_imag=16'b0010000001100101; end // in_theta = 0.831055 pi
 12'b011010100111: begin out_real=16'b1100100011000001; out_imag=16'b0010000001010000; end // in_theta = 0.831543 pi
 12'b011010101000: begin out_real=16'b1100100010110101; out_imag=16'b0010000000111010; end // in_theta = 0.832031 pi
 12'b011010101001: begin out_real=16'b1100100010101000; out_imag=16'b0010000000100100; end // in_theta = 0.832520 pi
 12'b011010101010: begin out_real=16'b1100100010011011; out_imag=16'b0010000000001111; end // in_theta = 0.833008 pi
 12'b011010101011: begin out_real=16'b1100100010001111; out_imag=16'b0001111111111001; end // in_theta = 0.833496 pi
 12'b011010101100: begin out_real=16'b1100100010000010; out_imag=16'b0001111111100011; end // in_theta = 0.833984 pi
 12'b011010101101: begin out_real=16'b1100100001110110; out_imag=16'b0001111111001101; end // in_theta = 0.834473 pi
 12'b011010101110: begin out_real=16'b1100100001101001; out_imag=16'b0001111110110111; end // in_theta = 0.834961 pi
 12'b011010101111: begin out_real=16'b1100100001011101; out_imag=16'b0001111110100010; end // in_theta = 0.835449 pi
 12'b011010110000: begin out_real=16'b1100100001010000; out_imag=16'b0001111110001100; end // in_theta = 0.835938 pi
 12'b011010110001: begin out_real=16'b1100100001000100; out_imag=16'b0001111101110110; end // in_theta = 0.836426 pi
 12'b011010110010: begin out_real=16'b1100100000111000; out_imag=16'b0001111101100000; end // in_theta = 0.836914 pi
 12'b011010110011: begin out_real=16'b1100100000101011; out_imag=16'b0001111101001010; end // in_theta = 0.837402 pi
 12'b011010110100: begin out_real=16'b1100100000011111; out_imag=16'b0001111100110100; end // in_theta = 0.837891 pi
 12'b011010110101: begin out_real=16'b1100100000010011; out_imag=16'b0001111100011110; end // in_theta = 0.838379 pi
 12'b011010110110: begin out_real=16'b1100100000000111; out_imag=16'b0001111100001000; end // in_theta = 0.838867 pi
 12'b011010110111: begin out_real=16'b1100011111111011; out_imag=16'b0001111011110010; end // in_theta = 0.839355 pi
 12'b011010111000: begin out_real=16'b1100011111101110; out_imag=16'b0001111011011100; end // in_theta = 0.839844 pi
 12'b011010111001: begin out_real=16'b1100011111100010; out_imag=16'b0001111011000110; end // in_theta = 0.840332 pi
 12'b011010111010: begin out_real=16'b1100011111010110; out_imag=16'b0001111010110000; end // in_theta = 0.840820 pi
 12'b011010111011: begin out_real=16'b1100011111001010; out_imag=16'b0001111010011010; end // in_theta = 0.841309 pi
 12'b011010111100: begin out_real=16'b1100011110111110; out_imag=16'b0001111010000100; end // in_theta = 0.841797 pi
 12'b011010111101: begin out_real=16'b1100011110110010; out_imag=16'b0001111001101110; end // in_theta = 0.842285 pi
 12'b011010111110: begin out_real=16'b1100011110100110; out_imag=16'b0001111001011000; end // in_theta = 0.842773 pi
 12'b011010111111: begin out_real=16'b1100011110011010; out_imag=16'b0001111001000010; end // in_theta = 0.843262 pi
 12'b011011000000: begin out_real=16'b1100011110001111; out_imag=16'b0001111000101011; end // in_theta = 0.843750 pi
 12'b011011000001: begin out_real=16'b1100011110000011; out_imag=16'b0001111000010101; end // in_theta = 0.844238 pi
 12'b011011000010: begin out_real=16'b1100011101110111; out_imag=16'b0001110111111111; end // in_theta = 0.844727 pi
 12'b011011000011: begin out_real=16'b1100011101101011; out_imag=16'b0001110111101001; end // in_theta = 0.845215 pi
 12'b011011000100: begin out_real=16'b1100011101011111; out_imag=16'b0001110111010011; end // in_theta = 0.845703 pi
 12'b011011000101: begin out_real=16'b1100011101010100; out_imag=16'b0001110110111100; end // in_theta = 0.846191 pi
 12'b011011000110: begin out_real=16'b1100011101001000; out_imag=16'b0001110110100110; end // in_theta = 0.846680 pi
 12'b011011000111: begin out_real=16'b1100011100111101; out_imag=16'b0001110110010000; end // in_theta = 0.847168 pi
 12'b011011001000: begin out_real=16'b1100011100110001; out_imag=16'b0001110101111001; end // in_theta = 0.847656 pi
 12'b011011001001: begin out_real=16'b1100011100100101; out_imag=16'b0001110101100011; end // in_theta = 0.848145 pi
 12'b011011001010: begin out_real=16'b1100011100011010; out_imag=16'b0001110101001101; end // in_theta = 0.848633 pi
 12'b011011001011: begin out_real=16'b1100011100001110; out_imag=16'b0001110100110110; end // in_theta = 0.849121 pi
 12'b011011001100: begin out_real=16'b1100011100000011; out_imag=16'b0001110100100000; end // in_theta = 0.849609 pi
 12'b011011001101: begin out_real=16'b1100011011110111; out_imag=16'b0001110100001010; end // in_theta = 0.850098 pi
 12'b011011001110: begin out_real=16'b1100011011101100; out_imag=16'b0001110011110011; end // in_theta = 0.850586 pi
 12'b011011001111: begin out_real=16'b1100011011100001; out_imag=16'b0001110011011101; end // in_theta = 0.851074 pi
 12'b011011010000: begin out_real=16'b1100011011010101; out_imag=16'b0001110011000110; end // in_theta = 0.851562 pi
 12'b011011010001: begin out_real=16'b1100011011001010; out_imag=16'b0001110010110000; end // in_theta = 0.852051 pi
 12'b011011010010: begin out_real=16'b1100011010111111; out_imag=16'b0001110010011001; end // in_theta = 0.852539 pi
 12'b011011010011: begin out_real=16'b1100011010110100; out_imag=16'b0001110010000011; end // in_theta = 0.853027 pi
 12'b011011010100: begin out_real=16'b1100011010101000; out_imag=16'b0001110001101100; end // in_theta = 0.853516 pi
 12'b011011010101: begin out_real=16'b1100011010011101; out_imag=16'b0001110001010110; end // in_theta = 0.854004 pi
 12'b011011010110: begin out_real=16'b1100011010010010; out_imag=16'b0001110000111111; end // in_theta = 0.854492 pi
 12'b011011010111: begin out_real=16'b1100011010000111; out_imag=16'b0001110000101001; end // in_theta = 0.854980 pi
 12'b011011011000: begin out_real=16'b1100011001111100; out_imag=16'b0001110000010010; end // in_theta = 0.855469 pi
 12'b011011011001: begin out_real=16'b1100011001110001; out_imag=16'b0001101111111100; end // in_theta = 0.855957 pi
 12'b011011011010: begin out_real=16'b1100011001100110; out_imag=16'b0001101111100101; end // in_theta = 0.856445 pi
 12'b011011011011: begin out_real=16'b1100011001011011; out_imag=16'b0001101111001110; end // in_theta = 0.856934 pi
 12'b011011011100: begin out_real=16'b1100011001010000; out_imag=16'b0001101110111000; end // in_theta = 0.857422 pi
 12'b011011011101: begin out_real=16'b1100011001000101; out_imag=16'b0001101110100001; end // in_theta = 0.857910 pi
 12'b011011011110: begin out_real=16'b1100011000111011; out_imag=16'b0001101110001010; end // in_theta = 0.858398 pi
 12'b011011011111: begin out_real=16'b1100011000110000; out_imag=16'b0001101101110100; end // in_theta = 0.858887 pi
 12'b011011100000: begin out_real=16'b1100011000100101; out_imag=16'b0001101101011101; end // in_theta = 0.859375 pi
 12'b011011100001: begin out_real=16'b1100011000011010; out_imag=16'b0001101101000110; end // in_theta = 0.859863 pi
 12'b011011100010: begin out_real=16'b1100011000010000; out_imag=16'b0001101100110000; end // in_theta = 0.860352 pi
 12'b011011100011: begin out_real=16'b1100011000000101; out_imag=16'b0001101100011001; end // in_theta = 0.860840 pi
 12'b011011100100: begin out_real=16'b1100010111111010; out_imag=16'b0001101100000010; end // in_theta = 0.861328 pi
 12'b011011100101: begin out_real=16'b1100010111110000; out_imag=16'b0001101011101011; end // in_theta = 0.861816 pi
 12'b011011100110: begin out_real=16'b1100010111100101; out_imag=16'b0001101011010100; end // in_theta = 0.862305 pi
 12'b011011100111: begin out_real=16'b1100010111011011; out_imag=16'b0001101010111110; end // in_theta = 0.862793 pi
 12'b011011101000: begin out_real=16'b1100010111010000; out_imag=16'b0001101010100111; end // in_theta = 0.863281 pi
 12'b011011101001: begin out_real=16'b1100010111000110; out_imag=16'b0001101010010000; end // in_theta = 0.863770 pi
 12'b011011101010: begin out_real=16'b1100010110111011; out_imag=16'b0001101001111001; end // in_theta = 0.864258 pi
 12'b011011101011: begin out_real=16'b1100010110110001; out_imag=16'b0001101001100010; end // in_theta = 0.864746 pi
 12'b011011101100: begin out_real=16'b1100010110100111; out_imag=16'b0001101001001011; end // in_theta = 0.865234 pi
 12'b011011101101: begin out_real=16'b1100010110011100; out_imag=16'b0001101000110100; end // in_theta = 0.865723 pi
 12'b011011101110: begin out_real=16'b1100010110010010; out_imag=16'b0001101000011101; end // in_theta = 0.866211 pi
 12'b011011101111: begin out_real=16'b1100010110001000; out_imag=16'b0001101000000110; end // in_theta = 0.866699 pi
 12'b011011110000: begin out_real=16'b1100010101111110; out_imag=16'b0001100111101111; end // in_theta = 0.867188 pi
 12'b011011110001: begin out_real=16'b1100010101110011; out_imag=16'b0001100111011000; end // in_theta = 0.867676 pi
 12'b011011110010: begin out_real=16'b1100010101101001; out_imag=16'b0001100111000001; end // in_theta = 0.868164 pi
 12'b011011110011: begin out_real=16'b1100010101011111; out_imag=16'b0001100110101010; end // in_theta = 0.868652 pi
 12'b011011110100: begin out_real=16'b1100010101010101; out_imag=16'b0001100110010011; end // in_theta = 0.869141 pi
 12'b011011110101: begin out_real=16'b1100010101001011; out_imag=16'b0001100101111100; end // in_theta = 0.869629 pi
 12'b011011110110: begin out_real=16'b1100010101000001; out_imag=16'b0001100101100101; end // in_theta = 0.870117 pi
 12'b011011110111: begin out_real=16'b1100010100110111; out_imag=16'b0001100101001110; end // in_theta = 0.870605 pi
 12'b011011111000: begin out_real=16'b1100010100101101; out_imag=16'b0001100100110111; end // in_theta = 0.871094 pi
 12'b011011111001: begin out_real=16'b1100010100100011; out_imag=16'b0001100100100000; end // in_theta = 0.871582 pi
 12'b011011111010: begin out_real=16'b1100010100011010; out_imag=16'b0001100100001001; end // in_theta = 0.872070 pi
 12'b011011111011: begin out_real=16'b1100010100010000; out_imag=16'b0001100011110010; end // in_theta = 0.872559 pi
 12'b011011111100: begin out_real=16'b1100010100000110; out_imag=16'b0001100011011011; end // in_theta = 0.873047 pi
 12'b011011111101: begin out_real=16'b1100010011111100; out_imag=16'b0001100011000011; end // in_theta = 0.873535 pi
 12'b011011111110: begin out_real=16'b1100010011110010; out_imag=16'b0001100010101100; end // in_theta = 0.874023 pi
 12'b011011111111: begin out_real=16'b1100010011101001; out_imag=16'b0001100010010101; end // in_theta = 0.874512 pi
 12'b011100000000: begin out_real=16'b1100010011011111; out_imag=16'b0001100001111110; end // in_theta = 0.875000 pi
 12'b011100000001: begin out_real=16'b1100010011010110; out_imag=16'b0001100001100111; end // in_theta = 0.875488 pi
 12'b011100000010: begin out_real=16'b1100010011001100; out_imag=16'b0001100001001111; end // in_theta = 0.875977 pi
 12'b011100000011: begin out_real=16'b1100010011000010; out_imag=16'b0001100000111000; end // in_theta = 0.876465 pi
 12'b011100000100: begin out_real=16'b1100010010111001; out_imag=16'b0001100000100001; end // in_theta = 0.876953 pi
 12'b011100000101: begin out_real=16'b1100010010110000; out_imag=16'b0001100000001010; end // in_theta = 0.877441 pi
 12'b011100000110: begin out_real=16'b1100010010100110; out_imag=16'b0001011111110010; end // in_theta = 0.877930 pi
 12'b011100000111: begin out_real=16'b1100010010011101; out_imag=16'b0001011111011011; end // in_theta = 0.878418 pi
 12'b011100001000: begin out_real=16'b1100010010010011; out_imag=16'b0001011111000100; end // in_theta = 0.878906 pi
 12'b011100001001: begin out_real=16'b1100010010001010; out_imag=16'b0001011110101100; end // in_theta = 0.879395 pi
 12'b011100001010: begin out_real=16'b1100010010000001; out_imag=16'b0001011110010101; end // in_theta = 0.879883 pi
 12'b011100001011: begin out_real=16'b1100010001111000; out_imag=16'b0001011101111110; end // in_theta = 0.880371 pi
 12'b011100001100: begin out_real=16'b1100010001101110; out_imag=16'b0001011101100110; end // in_theta = 0.880859 pi
 12'b011100001101: begin out_real=16'b1100010001100101; out_imag=16'b0001011101001111; end // in_theta = 0.881348 pi
 12'b011100001110: begin out_real=16'b1100010001011100; out_imag=16'b0001011100110111; end // in_theta = 0.881836 pi
 12'b011100001111: begin out_real=16'b1100010001010011; out_imag=16'b0001011100100000; end // in_theta = 0.882324 pi
 12'b011100010000: begin out_real=16'b1100010001001010; out_imag=16'b0001011100001001; end // in_theta = 0.882813 pi
 12'b011100010001: begin out_real=16'b1100010001000001; out_imag=16'b0001011011110001; end // in_theta = 0.883301 pi
 12'b011100010010: begin out_real=16'b1100010000111000; out_imag=16'b0001011011011010; end // in_theta = 0.883789 pi
 12'b011100010011: begin out_real=16'b1100010000101111; out_imag=16'b0001011011000010; end // in_theta = 0.884277 pi
 12'b011100010100: begin out_real=16'b1100010000100110; out_imag=16'b0001011010101011; end // in_theta = 0.884766 pi
 12'b011100010101: begin out_real=16'b1100010000011101; out_imag=16'b0001011010010011; end // in_theta = 0.885254 pi
 12'b011100010110: begin out_real=16'b1100010000010100; out_imag=16'b0001011001111100; end // in_theta = 0.885742 pi
 12'b011100010111: begin out_real=16'b1100010000001011; out_imag=16'b0001011001100100; end // in_theta = 0.886230 pi
 12'b011100011000: begin out_real=16'b1100010000000011; out_imag=16'b0001011001001100; end // in_theta = 0.886719 pi
 12'b011100011001: begin out_real=16'b1100001111111010; out_imag=16'b0001011000110101; end // in_theta = 0.887207 pi
 12'b011100011010: begin out_real=16'b1100001111110001; out_imag=16'b0001011000011101; end // in_theta = 0.887695 pi
 12'b011100011011: begin out_real=16'b1100001111101001; out_imag=16'b0001011000000110; end // in_theta = 0.888184 pi
 12'b011100011100: begin out_real=16'b1100001111100000; out_imag=16'b0001010111101110; end // in_theta = 0.888672 pi
 12'b011100011101: begin out_real=16'b1100001111010111; out_imag=16'b0001010111010111; end // in_theta = 0.889160 pi
 12'b011100011110: begin out_real=16'b1100001111001111; out_imag=16'b0001010110111111; end // in_theta = 0.889648 pi
 12'b011100011111: begin out_real=16'b1100001111000110; out_imag=16'b0001010110100111; end // in_theta = 0.890137 pi
 12'b011100100000: begin out_real=16'b1100001110111110; out_imag=16'b0001010110010000; end // in_theta = 0.890625 pi
 12'b011100100001: begin out_real=16'b1100001110110101; out_imag=16'b0001010101111000; end // in_theta = 0.891113 pi
 12'b011100100010: begin out_real=16'b1100001110101101; out_imag=16'b0001010101100000; end // in_theta = 0.891602 pi
 12'b011100100011: begin out_real=16'b1100001110100101; out_imag=16'b0001010101001001; end // in_theta = 0.892090 pi
 12'b011100100100: begin out_real=16'b1100001110011100; out_imag=16'b0001010100110001; end // in_theta = 0.892578 pi
 12'b011100100101: begin out_real=16'b1100001110010100; out_imag=16'b0001010100011001; end // in_theta = 0.893066 pi
 12'b011100100110: begin out_real=16'b1100001110001100; out_imag=16'b0001010100000001; end // in_theta = 0.893555 pi
 12'b011100100111: begin out_real=16'b1100001110000011; out_imag=16'b0001010011101010; end // in_theta = 0.894043 pi
 12'b011100101000: begin out_real=16'b1100001101111011; out_imag=16'b0001010011010010; end // in_theta = 0.894531 pi
 12'b011100101001: begin out_real=16'b1100001101110011; out_imag=16'b0001010010111010; end // in_theta = 0.895020 pi
 12'b011100101010: begin out_real=16'b1100001101101011; out_imag=16'b0001010010100010; end // in_theta = 0.895508 pi
 12'b011100101011: begin out_real=16'b1100001101100011; out_imag=16'b0001010010001011; end // in_theta = 0.895996 pi
 12'b011100101100: begin out_real=16'b1100001101011011; out_imag=16'b0001010001110011; end // in_theta = 0.896484 pi
 12'b011100101101: begin out_real=16'b1100001101010011; out_imag=16'b0001010001011011; end // in_theta = 0.896973 pi
 12'b011100101110: begin out_real=16'b1100001101001011; out_imag=16'b0001010001000011; end // in_theta = 0.897461 pi
 12'b011100101111: begin out_real=16'b1100001101000011; out_imag=16'b0001010000101011; end // in_theta = 0.897949 pi
 12'b011100110000: begin out_real=16'b1100001100111011; out_imag=16'b0001010000010011; end // in_theta = 0.898438 pi
 12'b011100110001: begin out_real=16'b1100001100110011; out_imag=16'b0001001111111011; end // in_theta = 0.898926 pi
 12'b011100110010: begin out_real=16'b1100001100101011; out_imag=16'b0001001111100100; end // in_theta = 0.899414 pi
 12'b011100110011: begin out_real=16'b1100001100100011; out_imag=16'b0001001111001100; end // in_theta = 0.899902 pi
 12'b011100110100: begin out_real=16'b1100001100011100; out_imag=16'b0001001110110100; end // in_theta = 0.900391 pi
 12'b011100110101: begin out_real=16'b1100001100010100; out_imag=16'b0001001110011100; end // in_theta = 0.900879 pi
 12'b011100110110: begin out_real=16'b1100001100001100; out_imag=16'b0001001110000100; end // in_theta = 0.901367 pi
 12'b011100110111: begin out_real=16'b1100001100000101; out_imag=16'b0001001101101100; end // in_theta = 0.901855 pi
 12'b011100111000: begin out_real=16'b1100001011111101; out_imag=16'b0001001101010100; end // in_theta = 0.902344 pi
 12'b011100111001: begin out_real=16'b1100001011110101; out_imag=16'b0001001100111100; end // in_theta = 0.902832 pi
 12'b011100111010: begin out_real=16'b1100001011101110; out_imag=16'b0001001100100100; end // in_theta = 0.903320 pi
 12'b011100111011: begin out_real=16'b1100001011100110; out_imag=16'b0001001100001100; end // in_theta = 0.903809 pi
 12'b011100111100: begin out_real=16'b1100001011011111; out_imag=16'b0001001011110100; end // in_theta = 0.904297 pi
 12'b011100111101: begin out_real=16'b1100001011011000; out_imag=16'b0001001011011100; end // in_theta = 0.904785 pi
 12'b011100111110: begin out_real=16'b1100001011010000; out_imag=16'b0001001011000100; end // in_theta = 0.905273 pi
 12'b011100111111: begin out_real=16'b1100001011001001; out_imag=16'b0001001010101100; end // in_theta = 0.905762 pi
 12'b011101000000: begin out_real=16'b1100001011000001; out_imag=16'b0001001010010100; end // in_theta = 0.906250 pi
 12'b011101000001: begin out_real=16'b1100001010111010; out_imag=16'b0001001001111100; end // in_theta = 0.906738 pi
 12'b011101000010: begin out_real=16'b1100001010110011; out_imag=16'b0001001001100100; end // in_theta = 0.907227 pi
 12'b011101000011: begin out_real=16'b1100001010101100; out_imag=16'b0001001001001100; end // in_theta = 0.907715 pi
 12'b011101000100: begin out_real=16'b1100001010100101; out_imag=16'b0001001000110100; end // in_theta = 0.908203 pi
 12'b011101000101: begin out_real=16'b1100001010011101; out_imag=16'b0001001000011100; end // in_theta = 0.908691 pi
 12'b011101000110: begin out_real=16'b1100001010010110; out_imag=16'b0001001000000100; end // in_theta = 0.909180 pi
 12'b011101000111: begin out_real=16'b1100001010001111; out_imag=16'b0001000111101011; end // in_theta = 0.909668 pi
 12'b011101001000: begin out_real=16'b1100001010001000; out_imag=16'b0001000111010011; end // in_theta = 0.910156 pi
 12'b011101001001: begin out_real=16'b1100001010000001; out_imag=16'b0001000110111011; end // in_theta = 0.910645 pi
 12'b011101001010: begin out_real=16'b1100001001111010; out_imag=16'b0001000110100011; end // in_theta = 0.911133 pi
 12'b011101001011: begin out_real=16'b1100001001110011; out_imag=16'b0001000110001011; end // in_theta = 0.911621 pi
 12'b011101001100: begin out_real=16'b1100001001101101; out_imag=16'b0001000101110011; end // in_theta = 0.912109 pi
 12'b011101001101: begin out_real=16'b1100001001100110; out_imag=16'b0001000101011010; end // in_theta = 0.912598 pi
 12'b011101001110: begin out_real=16'b1100001001011111; out_imag=16'b0001000101000010; end // in_theta = 0.913086 pi
 12'b011101001111: begin out_real=16'b1100001001011000; out_imag=16'b0001000100101010; end // in_theta = 0.913574 pi
 12'b011101010000: begin out_real=16'b1100001001010001; out_imag=16'b0001000100010010; end // in_theta = 0.914063 pi
 12'b011101010001: begin out_real=16'b1100001001001011; out_imag=16'b0001000011111010; end // in_theta = 0.914551 pi
 12'b011101010010: begin out_real=16'b1100001001000100; out_imag=16'b0001000011100001; end // in_theta = 0.915039 pi
 12'b011101010011: begin out_real=16'b1100001000111110; out_imag=16'b0001000011001001; end // in_theta = 0.915527 pi
 12'b011101010100: begin out_real=16'b1100001000110111; out_imag=16'b0001000010110001; end // in_theta = 0.916016 pi
 12'b011101010101: begin out_real=16'b1100001000110000; out_imag=16'b0001000010011001; end // in_theta = 0.916504 pi
 12'b011101010110: begin out_real=16'b1100001000101010; out_imag=16'b0001000010000000; end // in_theta = 0.916992 pi
 12'b011101010111: begin out_real=16'b1100001000100011; out_imag=16'b0001000001101000; end // in_theta = 0.917480 pi
 12'b011101011000: begin out_real=16'b1100001000011101; out_imag=16'b0001000001010000; end // in_theta = 0.917969 pi
 12'b011101011001: begin out_real=16'b1100001000010111; out_imag=16'b0001000000110111; end // in_theta = 0.918457 pi
 12'b011101011010: begin out_real=16'b1100001000010000; out_imag=16'b0001000000011111; end // in_theta = 0.918945 pi
 12'b011101011011: begin out_real=16'b1100001000001010; out_imag=16'b0001000000000111; end // in_theta = 0.919434 pi
 12'b011101011100: begin out_real=16'b1100001000000100; out_imag=16'b0000111111101110; end // in_theta = 0.919922 pi
 12'b011101011101: begin out_real=16'b1100000111111101; out_imag=16'b0000111111010110; end // in_theta = 0.920410 pi
 12'b011101011110: begin out_real=16'b1100000111110111; out_imag=16'b0000111110111110; end // in_theta = 0.920898 pi
 12'b011101011111: begin out_real=16'b1100000111110001; out_imag=16'b0000111110100101; end // in_theta = 0.921387 pi
 12'b011101100000: begin out_real=16'b1100000111101011; out_imag=16'b0000111110001101; end // in_theta = 0.921875 pi
 12'b011101100001: begin out_real=16'b1100000111100101; out_imag=16'b0000111101110101; end // in_theta = 0.922363 pi
 12'b011101100010: begin out_real=16'b1100000111011111; out_imag=16'b0000111101011100; end // in_theta = 0.922852 pi
 12'b011101100011: begin out_real=16'b1100000111011001; out_imag=16'b0000111101000100; end // in_theta = 0.923340 pi
 12'b011101100100: begin out_real=16'b1100000111010011; out_imag=16'b0000111100101011; end // in_theta = 0.923828 pi
 12'b011101100101: begin out_real=16'b1100000111001101; out_imag=16'b0000111100010011; end // in_theta = 0.924316 pi
 12'b011101100110: begin out_real=16'b1100000111000111; out_imag=16'b0000111011111011; end // in_theta = 0.924805 pi
 12'b011101100111: begin out_real=16'b1100000111000001; out_imag=16'b0000111011100010; end // in_theta = 0.925293 pi
 12'b011101101000: begin out_real=16'b1100000110111011; out_imag=16'b0000111011001010; end // in_theta = 0.925781 pi
 12'b011101101001: begin out_real=16'b1100000110110110; out_imag=16'b0000111010110001; end // in_theta = 0.926270 pi
 12'b011101101010: begin out_real=16'b1100000110110000; out_imag=16'b0000111010011001; end // in_theta = 0.926758 pi
 12'b011101101011: begin out_real=16'b1100000110101010; out_imag=16'b0000111010000000; end // in_theta = 0.927246 pi
 12'b011101101100: begin out_real=16'b1100000110100100; out_imag=16'b0000111001101000; end // in_theta = 0.927734 pi
 12'b011101101101: begin out_real=16'b1100000110011111; out_imag=16'b0000111001001111; end // in_theta = 0.928223 pi
 12'b011101101110: begin out_real=16'b1100000110011001; out_imag=16'b0000111000110111; end // in_theta = 0.928711 pi
 12'b011101101111: begin out_real=16'b1100000110010100; out_imag=16'b0000111000011110; end // in_theta = 0.929199 pi
 12'b011101110000: begin out_real=16'b1100000110001110; out_imag=16'b0000111000000110; end // in_theta = 0.929688 pi
 12'b011101110001: begin out_real=16'b1100000110001001; out_imag=16'b0000110111101101; end // in_theta = 0.930176 pi
 12'b011101110010: begin out_real=16'b1100000110000011; out_imag=16'b0000110111010101; end // in_theta = 0.930664 pi
 12'b011101110011: begin out_real=16'b1100000101111110; out_imag=16'b0000110110111100; end // in_theta = 0.931152 pi
 12'b011101110100: begin out_real=16'b1100000101111000; out_imag=16'b0000110110100100; end // in_theta = 0.931641 pi
 12'b011101110101: begin out_real=16'b1100000101110011; out_imag=16'b0000110110001011; end // in_theta = 0.932129 pi
 12'b011101110110: begin out_real=16'b1100000101101110; out_imag=16'b0000110101110010; end // in_theta = 0.932617 pi
 12'b011101110111: begin out_real=16'b1100000101101000; out_imag=16'b0000110101011010; end // in_theta = 0.933105 pi
 12'b011101111000: begin out_real=16'b1100000101100011; out_imag=16'b0000110101000001; end // in_theta = 0.933594 pi
 12'b011101111001: begin out_real=16'b1100000101011110; out_imag=16'b0000110100101001; end // in_theta = 0.934082 pi
 12'b011101111010: begin out_real=16'b1100000101011001; out_imag=16'b0000110100010000; end // in_theta = 0.934570 pi
 12'b011101111011: begin out_real=16'b1100000101010100; out_imag=16'b0000110011111000; end // in_theta = 0.935059 pi
 12'b011101111100: begin out_real=16'b1100000101001111; out_imag=16'b0000110011011111; end // in_theta = 0.935547 pi
 12'b011101111101: begin out_real=16'b1100000101001010; out_imag=16'b0000110011000110; end // in_theta = 0.936035 pi
 12'b011101111110: begin out_real=16'b1100000101000101; out_imag=16'b0000110010101110; end // in_theta = 0.936523 pi
 12'b011101111111: begin out_real=16'b1100000101000000; out_imag=16'b0000110010010101; end // in_theta = 0.937012 pi
 12'b011110000000: begin out_real=16'b1100000100111011; out_imag=16'b0000110001111100; end // in_theta = 0.937500 pi
 12'b011110000001: begin out_real=16'b1100000100110110; out_imag=16'b0000110001100100; end // in_theta = 0.937988 pi
 12'b011110000010: begin out_real=16'b1100000100110001; out_imag=16'b0000110001001011; end // in_theta = 0.938477 pi
 12'b011110000011: begin out_real=16'b1100000100101100; out_imag=16'b0000110000110010; end // in_theta = 0.938965 pi
 12'b011110000100: begin out_real=16'b1100000100101000; out_imag=16'b0000110000011010; end // in_theta = 0.939453 pi
 12'b011110000101: begin out_real=16'b1100000100100011; out_imag=16'b0000110000000001; end // in_theta = 0.939941 pi
 12'b011110000110: begin out_real=16'b1100000100011110; out_imag=16'b0000101111101000; end // in_theta = 0.940430 pi
 12'b011110000111: begin out_real=16'b1100000100011001; out_imag=16'b0000101111010000; end // in_theta = 0.940918 pi
 12'b011110001000: begin out_real=16'b1100000100010101; out_imag=16'b0000101110110111; end // in_theta = 0.941406 pi
 12'b011110001001: begin out_real=16'b1100000100010000; out_imag=16'b0000101110011110; end // in_theta = 0.941895 pi
 12'b011110001010: begin out_real=16'b1100000100001100; out_imag=16'b0000101110000101; end // in_theta = 0.942383 pi
 12'b011110001011: begin out_real=16'b1100000100000111; out_imag=16'b0000101101101101; end // in_theta = 0.942871 pi
 12'b011110001100: begin out_real=16'b1100000100000011; out_imag=16'b0000101101010100; end // in_theta = 0.943359 pi
 12'b011110001101: begin out_real=16'b1100000011111110; out_imag=16'b0000101100111011; end // in_theta = 0.943848 pi
 12'b011110001110: begin out_real=16'b1100000011111010; out_imag=16'b0000101100100011; end // in_theta = 0.944336 pi
 12'b011110001111: begin out_real=16'b1100000011110110; out_imag=16'b0000101100001010; end // in_theta = 0.944824 pi
 12'b011110010000: begin out_real=16'b1100000011110001; out_imag=16'b0000101011110001; end // in_theta = 0.945313 pi
 12'b011110010001: begin out_real=16'b1100000011101101; out_imag=16'b0000101011011000; end // in_theta = 0.945801 pi
 12'b011110010010: begin out_real=16'b1100000011101001; out_imag=16'b0000101011000000; end // in_theta = 0.946289 pi
 12'b011110010011: begin out_real=16'b1100000011100100; out_imag=16'b0000101010100111; end // in_theta = 0.946777 pi
 12'b011110010100: begin out_real=16'b1100000011100000; out_imag=16'b0000101010001110; end // in_theta = 0.947266 pi
 12'b011110010101: begin out_real=16'b1100000011011100; out_imag=16'b0000101001110101; end // in_theta = 0.947754 pi
 12'b011110010110: begin out_real=16'b1100000011011000; out_imag=16'b0000101001011100; end // in_theta = 0.948242 pi
 12'b011110010111: begin out_real=16'b1100000011010100; out_imag=16'b0000101001000100; end // in_theta = 0.948730 pi
 12'b011110011000: begin out_real=16'b1100000011010000; out_imag=16'b0000101000101011; end // in_theta = 0.949219 pi
 12'b011110011001: begin out_real=16'b1100000011001100; out_imag=16'b0000101000010010; end // in_theta = 0.949707 pi
 12'b011110011010: begin out_real=16'b1100000011001000; out_imag=16'b0000100111111001; end // in_theta = 0.950195 pi
 12'b011110011011: begin out_real=16'b1100000011000100; out_imag=16'b0000100111100000; end // in_theta = 0.950684 pi
 12'b011110011100: begin out_real=16'b1100000011000000; out_imag=16'b0000100111000111; end // in_theta = 0.951172 pi
 12'b011110011101: begin out_real=16'b1100000010111101; out_imag=16'b0000100110101111; end // in_theta = 0.951660 pi
 12'b011110011110: begin out_real=16'b1100000010111001; out_imag=16'b0000100110010110; end // in_theta = 0.952148 pi
 12'b011110011111: begin out_real=16'b1100000010110101; out_imag=16'b0000100101111101; end // in_theta = 0.952637 pi
 12'b011110100000: begin out_real=16'b1100000010110001; out_imag=16'b0000100101100100; end // in_theta = 0.953125 pi
 12'b011110100001: begin out_real=16'b1100000010101110; out_imag=16'b0000100101001011; end // in_theta = 0.953613 pi
 12'b011110100010: begin out_real=16'b1100000010101010; out_imag=16'b0000100100110010; end // in_theta = 0.954102 pi
 12'b011110100011: begin out_real=16'b1100000010100110; out_imag=16'b0000100100011001; end // in_theta = 0.954590 pi
 12'b011110100100: begin out_real=16'b1100000010100011; out_imag=16'b0000100100000001; end // in_theta = 0.955078 pi
 12'b011110100101: begin out_real=16'b1100000010011111; out_imag=16'b0000100011101000; end // in_theta = 0.955566 pi
 12'b011110100110: begin out_real=16'b1100000010011100; out_imag=16'b0000100011001111; end // in_theta = 0.956055 pi
 12'b011110100111: begin out_real=16'b1100000010011000; out_imag=16'b0000100010110110; end // in_theta = 0.956543 pi
 12'b011110101000: begin out_real=16'b1100000010010101; out_imag=16'b0000100010011101; end // in_theta = 0.957031 pi
 12'b011110101001: begin out_real=16'b1100000010010010; out_imag=16'b0000100010000100; end // in_theta = 0.957520 pi
 12'b011110101010: begin out_real=16'b1100000010001110; out_imag=16'b0000100001101011; end // in_theta = 0.958008 pi
 12'b011110101011: begin out_real=16'b1100000010001011; out_imag=16'b0000100001010010; end // in_theta = 0.958496 pi
 12'b011110101100: begin out_real=16'b1100000010001000; out_imag=16'b0000100000111001; end // in_theta = 0.958984 pi
 12'b011110101101: begin out_real=16'b1100000010000101; out_imag=16'b0000100000100000; end // in_theta = 0.959473 pi
 12'b011110101110: begin out_real=16'b1100000010000001; out_imag=16'b0000100000000111; end // in_theta = 0.959961 pi
 12'b011110101111: begin out_real=16'b1100000001111110; out_imag=16'b0000011111101111; end // in_theta = 0.960449 pi
 12'b011110110000: begin out_real=16'b1100000001111011; out_imag=16'b0000011111010110; end // in_theta = 0.960938 pi
 12'b011110110001: begin out_real=16'b1100000001111000; out_imag=16'b0000011110111101; end // in_theta = 0.961426 pi
 12'b011110110010: begin out_real=16'b1100000001110101; out_imag=16'b0000011110100100; end // in_theta = 0.961914 pi
 12'b011110110011: begin out_real=16'b1100000001110010; out_imag=16'b0000011110001011; end // in_theta = 0.962402 pi
 12'b011110110100: begin out_real=16'b1100000001101111; out_imag=16'b0000011101110010; end // in_theta = 0.962891 pi
 12'b011110110101: begin out_real=16'b1100000001101100; out_imag=16'b0000011101011001; end // in_theta = 0.963379 pi
 12'b011110110110: begin out_real=16'b1100000001101001; out_imag=16'b0000011101000000; end // in_theta = 0.963867 pi
 12'b011110110111: begin out_real=16'b1100000001100111; out_imag=16'b0000011100100111; end // in_theta = 0.964355 pi
 12'b011110111000: begin out_real=16'b1100000001100100; out_imag=16'b0000011100001110; end // in_theta = 0.964844 pi
 12'b011110111001: begin out_real=16'b1100000001100001; out_imag=16'b0000011011110101; end // in_theta = 0.965332 pi
 12'b011110111010: begin out_real=16'b1100000001011110; out_imag=16'b0000011011011100; end // in_theta = 0.965820 pi
 12'b011110111011: begin out_real=16'b1100000001011100; out_imag=16'b0000011011000011; end // in_theta = 0.966309 pi
 12'b011110111100: begin out_real=16'b1100000001011001; out_imag=16'b0000011010101010; end // in_theta = 0.966797 pi
 12'b011110111101: begin out_real=16'b1100000001010110; out_imag=16'b0000011010010001; end // in_theta = 0.967285 pi
 12'b011110111110: begin out_real=16'b1100000001010100; out_imag=16'b0000011001111000; end // in_theta = 0.967773 pi
 12'b011110111111: begin out_real=16'b1100000001010001; out_imag=16'b0000011001011111; end // in_theta = 0.968262 pi
 12'b011111000000: begin out_real=16'b1100000001001111; out_imag=16'b0000011001000110; end // in_theta = 0.968750 pi
 12'b011111000001: begin out_real=16'b1100000001001100; out_imag=16'b0000011000101101; end // in_theta = 0.969238 pi
 12'b011111000010: begin out_real=16'b1100000001001010; out_imag=16'b0000011000010100; end // in_theta = 0.969727 pi
 12'b011111000011: begin out_real=16'b1100000001001000; out_imag=16'b0000010111111011; end // in_theta = 0.970215 pi
 12'b011111000100: begin out_real=16'b1100000001000101; out_imag=16'b0000010111100010; end // in_theta = 0.970703 pi
 12'b011111000101: begin out_real=16'b1100000001000011; out_imag=16'b0000010111001001; end // in_theta = 0.971191 pi
 12'b011111000110: begin out_real=16'b1100000001000001; out_imag=16'b0000010110110000; end // in_theta = 0.971680 pi
 12'b011111000111: begin out_real=16'b1100000000111111; out_imag=16'b0000010110010111; end // in_theta = 0.972168 pi
 12'b011111001000: begin out_real=16'b1100000000111100; out_imag=16'b0000010101111110; end // in_theta = 0.972656 pi
 12'b011111001001: begin out_real=16'b1100000000111010; out_imag=16'b0000010101100101; end // in_theta = 0.973145 pi
 12'b011111001010: begin out_real=16'b1100000000111000; out_imag=16'b0000010101001100; end // in_theta = 0.973633 pi
 12'b011111001011: begin out_real=16'b1100000000110110; out_imag=16'b0000010100110011; end // in_theta = 0.974121 pi
 12'b011111001100: begin out_real=16'b1100000000110100; out_imag=16'b0000010100011010; end // in_theta = 0.974609 pi
 12'b011111001101: begin out_real=16'b1100000000110010; out_imag=16'b0000010100000000; end // in_theta = 0.975098 pi
 12'b011111001110: begin out_real=16'b1100000000110000; out_imag=16'b0000010011100111; end // in_theta = 0.975586 pi
 12'b011111001111: begin out_real=16'b1100000000101110; out_imag=16'b0000010011001110; end // in_theta = 0.976074 pi
 12'b011111010000: begin out_real=16'b1100000000101100; out_imag=16'b0000010010110101; end // in_theta = 0.976562 pi
 12'b011111010001: begin out_real=16'b1100000000101011; out_imag=16'b0000010010011100; end // in_theta = 0.977051 pi
 12'b011111010010: begin out_real=16'b1100000000101001; out_imag=16'b0000010010000011; end // in_theta = 0.977539 pi
 12'b011111010011: begin out_real=16'b1100000000100111; out_imag=16'b0000010001101010; end // in_theta = 0.978027 pi
 12'b011111010100: begin out_real=16'b1100000000100101; out_imag=16'b0000010001010001; end // in_theta = 0.978516 pi
 12'b011111010101: begin out_real=16'b1100000000100100; out_imag=16'b0000010000111000; end // in_theta = 0.979004 pi
 12'b011111010110: begin out_real=16'b1100000000100010; out_imag=16'b0000010000011111; end // in_theta = 0.979492 pi
 12'b011111010111: begin out_real=16'b1100000000100000; out_imag=16'b0000010000000110; end // in_theta = 0.979980 pi
 12'b011111011000: begin out_real=16'b1100000000011111; out_imag=16'b0000001111101101; end // in_theta = 0.980469 pi
 12'b011111011001: begin out_real=16'b1100000000011101; out_imag=16'b0000001111010100; end // in_theta = 0.980957 pi
 12'b011111011010: begin out_real=16'b1100000000011100; out_imag=16'b0000001110111011; end // in_theta = 0.981445 pi
 12'b011111011011: begin out_real=16'b1100000000011010; out_imag=16'b0000001110100001; end // in_theta = 0.981934 pi
 12'b011111011100: begin out_real=16'b1100000000011001; out_imag=16'b0000001110001000; end // in_theta = 0.982422 pi
 12'b011111011101: begin out_real=16'b1100000000011000; out_imag=16'b0000001101101111; end // in_theta = 0.982910 pi
 12'b011111011110: begin out_real=16'b1100000000010110; out_imag=16'b0000001101010110; end // in_theta = 0.983398 pi
 12'b011111011111: begin out_real=16'b1100000000010101; out_imag=16'b0000001100111101; end // in_theta = 0.983887 pi
 12'b011111100000: begin out_real=16'b1100000000010100; out_imag=16'b0000001100100100; end // in_theta = 0.984375 pi
 12'b011111100001: begin out_real=16'b1100000000010011; out_imag=16'b0000001100001011; end // in_theta = 0.984863 pi
 12'b011111100010: begin out_real=16'b1100000000010001; out_imag=16'b0000001011110010; end // in_theta = 0.985352 pi
 12'b011111100011: begin out_real=16'b1100000000010000; out_imag=16'b0000001011011001; end // in_theta = 0.985840 pi
 12'b011111100100: begin out_real=16'b1100000000001111; out_imag=16'b0000001011000000; end // in_theta = 0.986328 pi
 12'b011111100101: begin out_real=16'b1100000000001110; out_imag=16'b0000001010100110; end // in_theta = 0.986816 pi
 12'b011111100110: begin out_real=16'b1100000000001101; out_imag=16'b0000001010001101; end // in_theta = 0.987305 pi
 12'b011111100111: begin out_real=16'b1100000000001100; out_imag=16'b0000001001110100; end // in_theta = 0.987793 pi
 12'b011111101000: begin out_real=16'b1100000000001011; out_imag=16'b0000001001011011; end // in_theta = 0.988281 pi
 12'b011111101001: begin out_real=16'b1100000000001010; out_imag=16'b0000001001000010; end // in_theta = 0.988770 pi
 12'b011111101010: begin out_real=16'b1100000000001001; out_imag=16'b0000001000101001; end // in_theta = 0.989258 pi
 12'b011111101011: begin out_real=16'b1100000000001001; out_imag=16'b0000001000010000; end // in_theta = 0.989746 pi
 12'b011111101100: begin out_real=16'b1100000000001000; out_imag=16'b0000000111110111; end // in_theta = 0.990234 pi
 12'b011111101101: begin out_real=16'b1100000000000111; out_imag=16'b0000000111011101; end // in_theta = 0.990723 pi
 12'b011111101110: begin out_real=16'b1100000000000110; out_imag=16'b0000000111000100; end // in_theta = 0.991211 pi
 12'b011111101111: begin out_real=16'b1100000000000110; out_imag=16'b0000000110101011; end // in_theta = 0.991699 pi
 12'b011111110000: begin out_real=16'b1100000000000101; out_imag=16'b0000000110010010; end // in_theta = 0.992188 pi
 12'b011111110001: begin out_real=16'b1100000000000100; out_imag=16'b0000000101111001; end // in_theta = 0.992676 pi
 12'b011111110010: begin out_real=16'b1100000000000100; out_imag=16'b0000000101100000; end // in_theta = 0.993164 pi
 12'b011111110011: begin out_real=16'b1100000000000011; out_imag=16'b0000000101000111; end // in_theta = 0.993652 pi
 12'b011111110100: begin out_real=16'b1100000000000011; out_imag=16'b0000000100101110; end // in_theta = 0.994141 pi
 12'b011111110101: begin out_real=16'b1100000000000010; out_imag=16'b0000000100010100; end // in_theta = 0.994629 pi
 12'b011111110110: begin out_real=16'b1100000000000010; out_imag=16'b0000000011111011; end // in_theta = 0.995117 pi
 12'b011111110111: begin out_real=16'b1100000000000010; out_imag=16'b0000000011100010; end // in_theta = 0.995605 pi
 12'b011111111000: begin out_real=16'b1100000000000001; out_imag=16'b0000000011001001; end // in_theta = 0.996094 pi
 12'b011111111001: begin out_real=16'b1100000000000001; out_imag=16'b0000000010110000; end // in_theta = 0.996582 pi
 12'b011111111010: begin out_real=16'b1100000000000001; out_imag=16'b0000000010010111; end // in_theta = 0.997070 pi
 12'b011111111011: begin out_real=16'b1100000000000000; out_imag=16'b0000000001111110; end // in_theta = 0.997559 pi
 12'b011111111100: begin out_real=16'b1100000000000000; out_imag=16'b0000000001100101; end // in_theta = 0.998047 pi
 12'b011111111101: begin out_real=16'b1100000000000000; out_imag=16'b0000000001001011; end // in_theta = 0.998535 pi
 12'b011111111110: begin out_real=16'b1100000000000000; out_imag=16'b0000000000110010; end // in_theta = 0.999023 pi
 12'b011111111111: begin out_real=16'b1100000000000000; out_imag=16'b0000000000011001; end // in_theta = 0.999512 pi
 12'b100000000000: begin out_real=16'b1100000000000000; out_imag=16'b0000000000000000; end // in_theta = 1.000000 pi
 12'b100000000001: begin out_real=16'b1100000000000000; out_imag=16'b1111111111100111; end // in_theta = 1.000488 pi
 12'b100000000010: begin out_real=16'b1100000000000000; out_imag=16'b1111111111001110; end // in_theta = 1.000977 pi
 12'b100000000011: begin out_real=16'b1100000000000000; out_imag=16'b1111111110110101; end // in_theta = 1.001465 pi
 12'b100000000100: begin out_real=16'b1100000000000000; out_imag=16'b1111111110011011; end // in_theta = 1.001953 pi
 12'b100000000101: begin out_real=16'b1100000000000000; out_imag=16'b1111111110000010; end // in_theta = 1.002441 pi
 12'b100000000110: begin out_real=16'b1100000000000001; out_imag=16'b1111111101101001; end // in_theta = 1.002930 pi
 12'b100000000111: begin out_real=16'b1100000000000001; out_imag=16'b1111111101010000; end // in_theta = 1.003418 pi
 12'b100000001000: begin out_real=16'b1100000000000001; out_imag=16'b1111111100110111; end // in_theta = 1.003906 pi
 12'b100000001001: begin out_real=16'b1100000000000010; out_imag=16'b1111111100011110; end // in_theta = 1.004395 pi
 12'b100000001010: begin out_real=16'b1100000000000010; out_imag=16'b1111111100000101; end // in_theta = 1.004883 pi
 12'b100000001011: begin out_real=16'b1100000000000010; out_imag=16'b1111111011101100; end // in_theta = 1.005371 pi
 12'b100000001100: begin out_real=16'b1100000000000011; out_imag=16'b1111111011010010; end // in_theta = 1.005859 pi
 12'b100000001101: begin out_real=16'b1100000000000011; out_imag=16'b1111111010111001; end // in_theta = 1.006348 pi
 12'b100000001110: begin out_real=16'b1100000000000100; out_imag=16'b1111111010100000; end // in_theta = 1.006836 pi
 12'b100000001111: begin out_real=16'b1100000000000100; out_imag=16'b1111111010000111; end // in_theta = 1.007324 pi
 12'b100000010000: begin out_real=16'b1100000000000101; out_imag=16'b1111111001101110; end // in_theta = 1.007813 pi
 12'b100000010001: begin out_real=16'b1100000000000110; out_imag=16'b1111111001010101; end // in_theta = 1.008301 pi
 12'b100000010010: begin out_real=16'b1100000000000110; out_imag=16'b1111111000111100; end // in_theta = 1.008789 pi
 12'b100000010011: begin out_real=16'b1100000000000111; out_imag=16'b1111111000100011; end // in_theta = 1.009277 pi
 12'b100000010100: begin out_real=16'b1100000000001000; out_imag=16'b1111111000001001; end // in_theta = 1.009766 pi
 12'b100000010101: begin out_real=16'b1100000000001001; out_imag=16'b1111110111110000; end // in_theta = 1.010254 pi
 12'b100000010110: begin out_real=16'b1100000000001001; out_imag=16'b1111110111010111; end // in_theta = 1.010742 pi
 12'b100000010111: begin out_real=16'b1100000000001010; out_imag=16'b1111110110111110; end // in_theta = 1.011230 pi
 12'b100000011000: begin out_real=16'b1100000000001011; out_imag=16'b1111110110100101; end // in_theta = 1.011719 pi
 12'b100000011001: begin out_real=16'b1100000000001100; out_imag=16'b1111110110001100; end // in_theta = 1.012207 pi
 12'b100000011010: begin out_real=16'b1100000000001101; out_imag=16'b1111110101110011; end // in_theta = 1.012695 pi
 12'b100000011011: begin out_real=16'b1100000000001110; out_imag=16'b1111110101011010; end // in_theta = 1.013184 pi
 12'b100000011100: begin out_real=16'b1100000000001111; out_imag=16'b1111110101000000; end // in_theta = 1.013672 pi
 12'b100000011101: begin out_real=16'b1100000000010000; out_imag=16'b1111110100100111; end // in_theta = 1.014160 pi
 12'b100000011110: begin out_real=16'b1100000000010001; out_imag=16'b1111110100001110; end // in_theta = 1.014648 pi
 12'b100000011111: begin out_real=16'b1100000000010011; out_imag=16'b1111110011110101; end // in_theta = 1.015137 pi
 12'b100000100000: begin out_real=16'b1100000000010100; out_imag=16'b1111110011011100; end // in_theta = 1.015625 pi
 12'b100000100001: begin out_real=16'b1100000000010101; out_imag=16'b1111110011000011; end // in_theta = 1.016113 pi
 12'b100000100010: begin out_real=16'b1100000000010110; out_imag=16'b1111110010101010; end // in_theta = 1.016602 pi
 12'b100000100011: begin out_real=16'b1100000000011000; out_imag=16'b1111110010010001; end // in_theta = 1.017090 pi
 12'b100000100100: begin out_real=16'b1100000000011001; out_imag=16'b1111110001111000; end // in_theta = 1.017578 pi
 12'b100000100101: begin out_real=16'b1100000000011010; out_imag=16'b1111110001011111; end // in_theta = 1.018066 pi
 12'b100000100110: begin out_real=16'b1100000000011100; out_imag=16'b1111110001000101; end // in_theta = 1.018555 pi
 12'b100000100111: begin out_real=16'b1100000000011101; out_imag=16'b1111110000101100; end // in_theta = 1.019043 pi
 12'b100000101000: begin out_real=16'b1100000000011111; out_imag=16'b1111110000010011; end // in_theta = 1.019531 pi
 12'b100000101001: begin out_real=16'b1100000000100000; out_imag=16'b1111101111111010; end // in_theta = 1.020020 pi
 12'b100000101010: begin out_real=16'b1100000000100010; out_imag=16'b1111101111100001; end // in_theta = 1.020508 pi
 12'b100000101011: begin out_real=16'b1100000000100100; out_imag=16'b1111101111001000; end // in_theta = 1.020996 pi
 12'b100000101100: begin out_real=16'b1100000000100101; out_imag=16'b1111101110101111; end // in_theta = 1.021484 pi
 12'b100000101101: begin out_real=16'b1100000000100111; out_imag=16'b1111101110010110; end // in_theta = 1.021973 pi
 12'b100000101110: begin out_real=16'b1100000000101001; out_imag=16'b1111101101111101; end // in_theta = 1.022461 pi
 12'b100000101111: begin out_real=16'b1100000000101011; out_imag=16'b1111101101100100; end // in_theta = 1.022949 pi
 12'b100000110000: begin out_real=16'b1100000000101100; out_imag=16'b1111101101001011; end // in_theta = 1.023438 pi
 12'b100000110001: begin out_real=16'b1100000000101110; out_imag=16'b1111101100110010; end // in_theta = 1.023926 pi
 12'b100000110010: begin out_real=16'b1100000000110000; out_imag=16'b1111101100011001; end // in_theta = 1.024414 pi
 12'b100000110011: begin out_real=16'b1100000000110010; out_imag=16'b1111101100000000; end // in_theta = 1.024902 pi
 12'b100000110100: begin out_real=16'b1100000000110100; out_imag=16'b1111101011100110; end // in_theta = 1.025391 pi
 12'b100000110101: begin out_real=16'b1100000000110110; out_imag=16'b1111101011001101; end // in_theta = 1.025879 pi
 12'b100000110110: begin out_real=16'b1100000000111000; out_imag=16'b1111101010110100; end // in_theta = 1.026367 pi
 12'b100000110111: begin out_real=16'b1100000000111010; out_imag=16'b1111101010011011; end // in_theta = 1.026855 pi
 12'b100000111000: begin out_real=16'b1100000000111100; out_imag=16'b1111101010000010; end // in_theta = 1.027344 pi
 12'b100000111001: begin out_real=16'b1100000000111111; out_imag=16'b1111101001101001; end // in_theta = 1.027832 pi
 12'b100000111010: begin out_real=16'b1100000001000001; out_imag=16'b1111101001010000; end // in_theta = 1.028320 pi
 12'b100000111011: begin out_real=16'b1100000001000011; out_imag=16'b1111101000110111; end // in_theta = 1.028809 pi
 12'b100000111100: begin out_real=16'b1100000001000101; out_imag=16'b1111101000011110; end // in_theta = 1.029297 pi
 12'b100000111101: begin out_real=16'b1100000001001000; out_imag=16'b1111101000000101; end // in_theta = 1.029785 pi
 12'b100000111110: begin out_real=16'b1100000001001010; out_imag=16'b1111100111101100; end // in_theta = 1.030273 pi
 12'b100000111111: begin out_real=16'b1100000001001100; out_imag=16'b1111100111010011; end // in_theta = 1.030762 pi
 12'b100001000000: begin out_real=16'b1100000001001111; out_imag=16'b1111100110111010; end // in_theta = 1.031250 pi
 12'b100001000001: begin out_real=16'b1100000001010001; out_imag=16'b1111100110100001; end // in_theta = 1.031738 pi
 12'b100001000010: begin out_real=16'b1100000001010100; out_imag=16'b1111100110001000; end // in_theta = 1.032227 pi
 12'b100001000011: begin out_real=16'b1100000001010110; out_imag=16'b1111100101101111; end // in_theta = 1.032715 pi
 12'b100001000100: begin out_real=16'b1100000001011001; out_imag=16'b1111100101010110; end // in_theta = 1.033203 pi
 12'b100001000101: begin out_real=16'b1100000001011100; out_imag=16'b1111100100111101; end // in_theta = 1.033691 pi
 12'b100001000110: begin out_real=16'b1100000001011110; out_imag=16'b1111100100100100; end // in_theta = 1.034180 pi
 12'b100001000111: begin out_real=16'b1100000001100001; out_imag=16'b1111100100001011; end // in_theta = 1.034668 pi
 12'b100001001000: begin out_real=16'b1100000001100100; out_imag=16'b1111100011110010; end // in_theta = 1.035156 pi
 12'b100001001001: begin out_real=16'b1100000001100111; out_imag=16'b1111100011011001; end // in_theta = 1.035645 pi
 12'b100001001010: begin out_real=16'b1100000001101001; out_imag=16'b1111100011000000; end // in_theta = 1.036133 pi
 12'b100001001011: begin out_real=16'b1100000001101100; out_imag=16'b1111100010100111; end // in_theta = 1.036621 pi
 12'b100001001100: begin out_real=16'b1100000001101111; out_imag=16'b1111100010001110; end // in_theta = 1.037109 pi
 12'b100001001101: begin out_real=16'b1100000001110010; out_imag=16'b1111100001110101; end // in_theta = 1.037598 pi
 12'b100001001110: begin out_real=16'b1100000001110101; out_imag=16'b1111100001011100; end // in_theta = 1.038086 pi
 12'b100001001111: begin out_real=16'b1100000001111000; out_imag=16'b1111100001000011; end // in_theta = 1.038574 pi
 12'b100001010000: begin out_real=16'b1100000001111011; out_imag=16'b1111100000101010; end // in_theta = 1.039063 pi
 12'b100001010001: begin out_real=16'b1100000001111110; out_imag=16'b1111100000010001; end // in_theta = 1.039551 pi
 12'b100001010010: begin out_real=16'b1100000010000001; out_imag=16'b1111011111111001; end // in_theta = 1.040039 pi
 12'b100001010011: begin out_real=16'b1100000010000101; out_imag=16'b1111011111100000; end // in_theta = 1.040527 pi
 12'b100001010100: begin out_real=16'b1100000010001000; out_imag=16'b1111011111000111; end // in_theta = 1.041016 pi
 12'b100001010101: begin out_real=16'b1100000010001011; out_imag=16'b1111011110101110; end // in_theta = 1.041504 pi
 12'b100001010110: begin out_real=16'b1100000010001110; out_imag=16'b1111011110010101; end // in_theta = 1.041992 pi
 12'b100001010111: begin out_real=16'b1100000010010010; out_imag=16'b1111011101111100; end // in_theta = 1.042480 pi
 12'b100001011000: begin out_real=16'b1100000010010101; out_imag=16'b1111011101100011; end // in_theta = 1.042969 pi
 12'b100001011001: begin out_real=16'b1100000010011000; out_imag=16'b1111011101001010; end // in_theta = 1.043457 pi
 12'b100001011010: begin out_real=16'b1100000010011100; out_imag=16'b1111011100110001; end // in_theta = 1.043945 pi
 12'b100001011011: begin out_real=16'b1100000010011111; out_imag=16'b1111011100011000; end // in_theta = 1.044434 pi
 12'b100001011100: begin out_real=16'b1100000010100011; out_imag=16'b1111011011111111; end // in_theta = 1.044922 pi
 12'b100001011101: begin out_real=16'b1100000010100110; out_imag=16'b1111011011100111; end // in_theta = 1.045410 pi
 12'b100001011110: begin out_real=16'b1100000010101010; out_imag=16'b1111011011001110; end // in_theta = 1.045898 pi
 12'b100001011111: begin out_real=16'b1100000010101110; out_imag=16'b1111011010110101; end // in_theta = 1.046387 pi
 12'b100001100000: begin out_real=16'b1100000010110001; out_imag=16'b1111011010011100; end // in_theta = 1.046875 pi
 12'b100001100001: begin out_real=16'b1100000010110101; out_imag=16'b1111011010000011; end // in_theta = 1.047363 pi
 12'b100001100010: begin out_real=16'b1100000010111001; out_imag=16'b1111011001101010; end // in_theta = 1.047852 pi
 12'b100001100011: begin out_real=16'b1100000010111101; out_imag=16'b1111011001010001; end // in_theta = 1.048340 pi
 12'b100001100100: begin out_real=16'b1100000011000000; out_imag=16'b1111011000111001; end // in_theta = 1.048828 pi
 12'b100001100101: begin out_real=16'b1100000011000100; out_imag=16'b1111011000100000; end // in_theta = 1.049316 pi
 12'b100001100110: begin out_real=16'b1100000011001000; out_imag=16'b1111011000000111; end // in_theta = 1.049805 pi
 12'b100001100111: begin out_real=16'b1100000011001100; out_imag=16'b1111010111101110; end // in_theta = 1.050293 pi
 12'b100001101000: begin out_real=16'b1100000011010000; out_imag=16'b1111010111010101; end // in_theta = 1.050781 pi
 12'b100001101001: begin out_real=16'b1100000011010100; out_imag=16'b1111010110111100; end // in_theta = 1.051270 pi
 12'b100001101010: begin out_real=16'b1100000011011000; out_imag=16'b1111010110100100; end // in_theta = 1.051758 pi
 12'b100001101011: begin out_real=16'b1100000011011100; out_imag=16'b1111010110001011; end // in_theta = 1.052246 pi
 12'b100001101100: begin out_real=16'b1100000011100000; out_imag=16'b1111010101110010; end // in_theta = 1.052734 pi
 12'b100001101101: begin out_real=16'b1100000011100100; out_imag=16'b1111010101011001; end // in_theta = 1.053223 pi
 12'b100001101110: begin out_real=16'b1100000011101001; out_imag=16'b1111010101000000; end // in_theta = 1.053711 pi
 12'b100001101111: begin out_real=16'b1100000011101101; out_imag=16'b1111010100101000; end // in_theta = 1.054199 pi
 12'b100001110000: begin out_real=16'b1100000011110001; out_imag=16'b1111010100001111; end // in_theta = 1.054688 pi
 12'b100001110001: begin out_real=16'b1100000011110110; out_imag=16'b1111010011110110; end // in_theta = 1.055176 pi
 12'b100001110010: begin out_real=16'b1100000011111010; out_imag=16'b1111010011011101; end // in_theta = 1.055664 pi
 12'b100001110011: begin out_real=16'b1100000011111110; out_imag=16'b1111010011000101; end // in_theta = 1.056152 pi
 12'b100001110100: begin out_real=16'b1100000100000011; out_imag=16'b1111010010101100; end // in_theta = 1.056641 pi
 12'b100001110101: begin out_real=16'b1100000100000111; out_imag=16'b1111010010010011; end // in_theta = 1.057129 pi
 12'b100001110110: begin out_real=16'b1100000100001100; out_imag=16'b1111010001111011; end // in_theta = 1.057617 pi
 12'b100001110111: begin out_real=16'b1100000100010000; out_imag=16'b1111010001100010; end // in_theta = 1.058105 pi
 12'b100001111000: begin out_real=16'b1100000100010101; out_imag=16'b1111010001001001; end // in_theta = 1.058594 pi
 12'b100001111001: begin out_real=16'b1100000100011001; out_imag=16'b1111010000110000; end // in_theta = 1.059082 pi
 12'b100001111010: begin out_real=16'b1100000100011110; out_imag=16'b1111010000011000; end // in_theta = 1.059570 pi
 12'b100001111011: begin out_real=16'b1100000100100011; out_imag=16'b1111001111111111; end // in_theta = 1.060059 pi
 12'b100001111100: begin out_real=16'b1100000100101000; out_imag=16'b1111001111100110; end // in_theta = 1.060547 pi
 12'b100001111101: begin out_real=16'b1100000100101100; out_imag=16'b1111001111001110; end // in_theta = 1.061035 pi
 12'b100001111110: begin out_real=16'b1100000100110001; out_imag=16'b1111001110110101; end // in_theta = 1.061523 pi
 12'b100001111111: begin out_real=16'b1100000100110110; out_imag=16'b1111001110011100; end // in_theta = 1.062012 pi
 12'b100010000000: begin out_real=16'b1100000100111011; out_imag=16'b1111001110000100; end // in_theta = 1.062500 pi
 12'b100010000001: begin out_real=16'b1100000101000000; out_imag=16'b1111001101101011; end // in_theta = 1.062988 pi
 12'b100010000010: begin out_real=16'b1100000101000101; out_imag=16'b1111001101010010; end // in_theta = 1.063477 pi
 12'b100010000011: begin out_real=16'b1100000101001010; out_imag=16'b1111001100111010; end // in_theta = 1.063965 pi
 12'b100010000100: begin out_real=16'b1100000101001111; out_imag=16'b1111001100100001; end // in_theta = 1.064453 pi
 12'b100010000101: begin out_real=16'b1100000101010100; out_imag=16'b1111001100001000; end // in_theta = 1.064941 pi
 12'b100010000110: begin out_real=16'b1100000101011001; out_imag=16'b1111001011110000; end // in_theta = 1.065430 pi
 12'b100010000111: begin out_real=16'b1100000101011110; out_imag=16'b1111001011010111; end // in_theta = 1.065918 pi
 12'b100010001000: begin out_real=16'b1100000101100011; out_imag=16'b1111001010111111; end // in_theta = 1.066406 pi
 12'b100010001001: begin out_real=16'b1100000101101000; out_imag=16'b1111001010100110; end // in_theta = 1.066895 pi
 12'b100010001010: begin out_real=16'b1100000101101110; out_imag=16'b1111001010001110; end // in_theta = 1.067383 pi
 12'b100010001011: begin out_real=16'b1100000101110011; out_imag=16'b1111001001110101; end // in_theta = 1.067871 pi
 12'b100010001100: begin out_real=16'b1100000101111000; out_imag=16'b1111001001011100; end // in_theta = 1.068359 pi
 12'b100010001101: begin out_real=16'b1100000101111110; out_imag=16'b1111001001000100; end // in_theta = 1.068848 pi
 12'b100010001110: begin out_real=16'b1100000110000011; out_imag=16'b1111001000101011; end // in_theta = 1.069336 pi
 12'b100010001111: begin out_real=16'b1100000110001001; out_imag=16'b1111001000010011; end // in_theta = 1.069824 pi
 12'b100010010000: begin out_real=16'b1100000110001110; out_imag=16'b1111000111111010; end // in_theta = 1.070313 pi
 12'b100010010001: begin out_real=16'b1100000110010100; out_imag=16'b1111000111100010; end // in_theta = 1.070801 pi
 12'b100010010010: begin out_real=16'b1100000110011001; out_imag=16'b1111000111001001; end // in_theta = 1.071289 pi
 12'b100010010011: begin out_real=16'b1100000110011111; out_imag=16'b1111000110110001; end // in_theta = 1.071777 pi
 12'b100010010100: begin out_real=16'b1100000110100100; out_imag=16'b1111000110011000; end // in_theta = 1.072266 pi
 12'b100010010101: begin out_real=16'b1100000110101010; out_imag=16'b1111000110000000; end // in_theta = 1.072754 pi
 12'b100010010110: begin out_real=16'b1100000110110000; out_imag=16'b1111000101100111; end // in_theta = 1.073242 pi
 12'b100010010111: begin out_real=16'b1100000110110110; out_imag=16'b1111000101001111; end // in_theta = 1.073730 pi
 12'b100010011000: begin out_real=16'b1100000110111011; out_imag=16'b1111000100110110; end // in_theta = 1.074219 pi
 12'b100010011001: begin out_real=16'b1100000111000001; out_imag=16'b1111000100011110; end // in_theta = 1.074707 pi
 12'b100010011010: begin out_real=16'b1100000111000111; out_imag=16'b1111000100000101; end // in_theta = 1.075195 pi
 12'b100010011011: begin out_real=16'b1100000111001101; out_imag=16'b1111000011101101; end // in_theta = 1.075684 pi
 12'b100010011100: begin out_real=16'b1100000111010011; out_imag=16'b1111000011010101; end // in_theta = 1.076172 pi
 12'b100010011101: begin out_real=16'b1100000111011001; out_imag=16'b1111000010111100; end // in_theta = 1.076660 pi
 12'b100010011110: begin out_real=16'b1100000111011111; out_imag=16'b1111000010100100; end // in_theta = 1.077148 pi
 12'b100010011111: begin out_real=16'b1100000111100101; out_imag=16'b1111000010001011; end // in_theta = 1.077637 pi
 12'b100010100000: begin out_real=16'b1100000111101011; out_imag=16'b1111000001110011; end // in_theta = 1.078125 pi
 12'b100010100001: begin out_real=16'b1100000111110001; out_imag=16'b1111000001011011; end // in_theta = 1.078613 pi
 12'b100010100010: begin out_real=16'b1100000111110111; out_imag=16'b1111000001000010; end // in_theta = 1.079102 pi
 12'b100010100011: begin out_real=16'b1100000111111101; out_imag=16'b1111000000101010; end // in_theta = 1.079590 pi
 12'b100010100100: begin out_real=16'b1100001000000100; out_imag=16'b1111000000010010; end // in_theta = 1.080078 pi
 12'b100010100101: begin out_real=16'b1100001000001010; out_imag=16'b1110111111111001; end // in_theta = 1.080566 pi
 12'b100010100110: begin out_real=16'b1100001000010000; out_imag=16'b1110111111100001; end // in_theta = 1.081055 pi
 12'b100010100111: begin out_real=16'b1100001000010111; out_imag=16'b1110111111001001; end // in_theta = 1.081543 pi
 12'b100010101000: begin out_real=16'b1100001000011101; out_imag=16'b1110111110110000; end // in_theta = 1.082031 pi
 12'b100010101001: begin out_real=16'b1100001000100011; out_imag=16'b1110111110011000; end // in_theta = 1.082520 pi
 12'b100010101010: begin out_real=16'b1100001000101010; out_imag=16'b1110111110000000; end // in_theta = 1.083008 pi
 12'b100010101011: begin out_real=16'b1100001000110000; out_imag=16'b1110111101100111; end // in_theta = 1.083496 pi
 12'b100010101100: begin out_real=16'b1100001000110111; out_imag=16'b1110111101001111; end // in_theta = 1.083984 pi
 12'b100010101101: begin out_real=16'b1100001000111110; out_imag=16'b1110111100110111; end // in_theta = 1.084473 pi
 12'b100010101110: begin out_real=16'b1100001001000100; out_imag=16'b1110111100011111; end // in_theta = 1.084961 pi
 12'b100010101111: begin out_real=16'b1100001001001011; out_imag=16'b1110111100000110; end // in_theta = 1.085449 pi
 12'b100010110000: begin out_real=16'b1100001001010001; out_imag=16'b1110111011101110; end // in_theta = 1.085938 pi
 12'b100010110001: begin out_real=16'b1100001001011000; out_imag=16'b1110111011010110; end // in_theta = 1.086426 pi
 12'b100010110010: begin out_real=16'b1100001001011111; out_imag=16'b1110111010111110; end // in_theta = 1.086914 pi
 12'b100010110011: begin out_real=16'b1100001001100110; out_imag=16'b1110111010100110; end // in_theta = 1.087402 pi
 12'b100010110100: begin out_real=16'b1100001001101101; out_imag=16'b1110111010001101; end // in_theta = 1.087891 pi
 12'b100010110101: begin out_real=16'b1100001001110011; out_imag=16'b1110111001110101; end // in_theta = 1.088379 pi
 12'b100010110110: begin out_real=16'b1100001001111010; out_imag=16'b1110111001011101; end // in_theta = 1.088867 pi
 12'b100010110111: begin out_real=16'b1100001010000001; out_imag=16'b1110111001000101; end // in_theta = 1.089355 pi
 12'b100010111000: begin out_real=16'b1100001010001000; out_imag=16'b1110111000101101; end // in_theta = 1.089844 pi
 12'b100010111001: begin out_real=16'b1100001010001111; out_imag=16'b1110111000010101; end // in_theta = 1.090332 pi
 12'b100010111010: begin out_real=16'b1100001010010110; out_imag=16'b1110110111111100; end // in_theta = 1.090820 pi
 12'b100010111011: begin out_real=16'b1100001010011101; out_imag=16'b1110110111100100; end // in_theta = 1.091309 pi
 12'b100010111100: begin out_real=16'b1100001010100101; out_imag=16'b1110110111001100; end // in_theta = 1.091797 pi
 12'b100010111101: begin out_real=16'b1100001010101100; out_imag=16'b1110110110110100; end // in_theta = 1.092285 pi
 12'b100010111110: begin out_real=16'b1100001010110011; out_imag=16'b1110110110011100; end // in_theta = 1.092773 pi
 12'b100010111111: begin out_real=16'b1100001010111010; out_imag=16'b1110110110000100; end // in_theta = 1.093262 pi
 12'b100011000000: begin out_real=16'b1100001011000001; out_imag=16'b1110110101101100; end // in_theta = 1.093750 pi
 12'b100011000001: begin out_real=16'b1100001011001001; out_imag=16'b1110110101010100; end // in_theta = 1.094238 pi
 12'b100011000010: begin out_real=16'b1100001011010000; out_imag=16'b1110110100111100; end // in_theta = 1.094727 pi
 12'b100011000011: begin out_real=16'b1100001011011000; out_imag=16'b1110110100100100; end // in_theta = 1.095215 pi
 12'b100011000100: begin out_real=16'b1100001011011111; out_imag=16'b1110110100001100; end // in_theta = 1.095703 pi
 12'b100011000101: begin out_real=16'b1100001011100110; out_imag=16'b1110110011110100; end // in_theta = 1.096191 pi
 12'b100011000110: begin out_real=16'b1100001011101110; out_imag=16'b1110110011011100; end // in_theta = 1.096680 pi
 12'b100011000111: begin out_real=16'b1100001011110101; out_imag=16'b1110110011000100; end // in_theta = 1.097168 pi
 12'b100011001000: begin out_real=16'b1100001011111101; out_imag=16'b1110110010101100; end // in_theta = 1.097656 pi
 12'b100011001001: begin out_real=16'b1100001100000101; out_imag=16'b1110110010010100; end // in_theta = 1.098145 pi
 12'b100011001010: begin out_real=16'b1100001100001100; out_imag=16'b1110110001111100; end // in_theta = 1.098633 pi
 12'b100011001011: begin out_real=16'b1100001100010100; out_imag=16'b1110110001100100; end // in_theta = 1.099121 pi
 12'b100011001100: begin out_real=16'b1100001100011100; out_imag=16'b1110110001001100; end // in_theta = 1.099609 pi
 12'b100011001101: begin out_real=16'b1100001100100011; out_imag=16'b1110110000110100; end // in_theta = 1.100098 pi
 12'b100011001110: begin out_real=16'b1100001100101011; out_imag=16'b1110110000011100; end // in_theta = 1.100586 pi
 12'b100011001111: begin out_real=16'b1100001100110011; out_imag=16'b1110110000000101; end // in_theta = 1.101074 pi
 12'b100011010000: begin out_real=16'b1100001100111011; out_imag=16'b1110101111101101; end // in_theta = 1.101563 pi
 12'b100011010001: begin out_real=16'b1100001101000011; out_imag=16'b1110101111010101; end // in_theta = 1.102051 pi
 12'b100011010010: begin out_real=16'b1100001101001011; out_imag=16'b1110101110111101; end // in_theta = 1.102539 pi
 12'b100011010011: begin out_real=16'b1100001101010011; out_imag=16'b1110101110100101; end // in_theta = 1.103027 pi
 12'b100011010100: begin out_real=16'b1100001101011011; out_imag=16'b1110101110001101; end // in_theta = 1.103516 pi
 12'b100011010101: begin out_real=16'b1100001101100011; out_imag=16'b1110101101110101; end // in_theta = 1.104004 pi
 12'b100011010110: begin out_real=16'b1100001101101011; out_imag=16'b1110101101011110; end // in_theta = 1.104492 pi
 12'b100011010111: begin out_real=16'b1100001101110011; out_imag=16'b1110101101000110; end // in_theta = 1.104980 pi
 12'b100011011000: begin out_real=16'b1100001101111011; out_imag=16'b1110101100101110; end // in_theta = 1.105469 pi
 12'b100011011001: begin out_real=16'b1100001110000011; out_imag=16'b1110101100010110; end // in_theta = 1.105957 pi
 12'b100011011010: begin out_real=16'b1100001110001100; out_imag=16'b1110101011111111; end // in_theta = 1.106445 pi
 12'b100011011011: begin out_real=16'b1100001110010100; out_imag=16'b1110101011100111; end // in_theta = 1.106934 pi
 12'b100011011100: begin out_real=16'b1100001110011100; out_imag=16'b1110101011001111; end // in_theta = 1.107422 pi
 12'b100011011101: begin out_real=16'b1100001110100101; out_imag=16'b1110101010110111; end // in_theta = 1.107910 pi
 12'b100011011110: begin out_real=16'b1100001110101101; out_imag=16'b1110101010100000; end // in_theta = 1.108398 pi
 12'b100011011111: begin out_real=16'b1100001110110101; out_imag=16'b1110101010001000; end // in_theta = 1.108887 pi
 12'b100011100000: begin out_real=16'b1100001110111110; out_imag=16'b1110101001110000; end // in_theta = 1.109375 pi
 12'b100011100001: begin out_real=16'b1100001111000110; out_imag=16'b1110101001011001; end // in_theta = 1.109863 pi
 12'b100011100010: begin out_real=16'b1100001111001111; out_imag=16'b1110101001000001; end // in_theta = 1.110352 pi
 12'b100011100011: begin out_real=16'b1100001111010111; out_imag=16'b1110101000101001; end // in_theta = 1.110840 pi
 12'b100011100100: begin out_real=16'b1100001111100000; out_imag=16'b1110101000010010; end // in_theta = 1.111328 pi
 12'b100011100101: begin out_real=16'b1100001111101001; out_imag=16'b1110100111111010; end // in_theta = 1.111816 pi
 12'b100011100110: begin out_real=16'b1100001111110001; out_imag=16'b1110100111100011; end // in_theta = 1.112305 pi
 12'b100011100111: begin out_real=16'b1100001111111010; out_imag=16'b1110100111001011; end // in_theta = 1.112793 pi
 12'b100011101000: begin out_real=16'b1100010000000011; out_imag=16'b1110100110110100; end // in_theta = 1.113281 pi
 12'b100011101001: begin out_real=16'b1100010000001011; out_imag=16'b1110100110011100; end // in_theta = 1.113770 pi
 12'b100011101010: begin out_real=16'b1100010000010100; out_imag=16'b1110100110000100; end // in_theta = 1.114258 pi
 12'b100011101011: begin out_real=16'b1100010000011101; out_imag=16'b1110100101101101; end // in_theta = 1.114746 pi
 12'b100011101100: begin out_real=16'b1100010000100110; out_imag=16'b1110100101010101; end // in_theta = 1.115234 pi
 12'b100011101101: begin out_real=16'b1100010000101111; out_imag=16'b1110100100111110; end // in_theta = 1.115723 pi
 12'b100011101110: begin out_real=16'b1100010000111000; out_imag=16'b1110100100100110; end // in_theta = 1.116211 pi
 12'b100011101111: begin out_real=16'b1100010001000001; out_imag=16'b1110100100001111; end // in_theta = 1.116699 pi
 12'b100011110000: begin out_real=16'b1100010001001010; out_imag=16'b1110100011110111; end // in_theta = 1.117188 pi
 12'b100011110001: begin out_real=16'b1100010001010011; out_imag=16'b1110100011100000; end // in_theta = 1.117676 pi
 12'b100011110010: begin out_real=16'b1100010001011100; out_imag=16'b1110100011001001; end // in_theta = 1.118164 pi
 12'b100011110011: begin out_real=16'b1100010001100101; out_imag=16'b1110100010110001; end // in_theta = 1.118652 pi
 12'b100011110100: begin out_real=16'b1100010001101110; out_imag=16'b1110100010011010; end // in_theta = 1.119141 pi
 12'b100011110101: begin out_real=16'b1100010001111000; out_imag=16'b1110100010000010; end // in_theta = 1.119629 pi
 12'b100011110110: begin out_real=16'b1100010010000001; out_imag=16'b1110100001101011; end // in_theta = 1.120117 pi
 12'b100011110111: begin out_real=16'b1100010010001010; out_imag=16'b1110100001010100; end // in_theta = 1.120605 pi
 12'b100011111000: begin out_real=16'b1100010010010011; out_imag=16'b1110100000111100; end // in_theta = 1.121094 pi
 12'b100011111001: begin out_real=16'b1100010010011101; out_imag=16'b1110100000100101; end // in_theta = 1.121582 pi
 12'b100011111010: begin out_real=16'b1100010010100110; out_imag=16'b1110100000001110; end // in_theta = 1.122070 pi
 12'b100011111011: begin out_real=16'b1100010010110000; out_imag=16'b1110011111110110; end // in_theta = 1.122559 pi
 12'b100011111100: begin out_real=16'b1100010010111001; out_imag=16'b1110011111011111; end // in_theta = 1.123047 pi
 12'b100011111101: begin out_real=16'b1100010011000010; out_imag=16'b1110011111001000; end // in_theta = 1.123535 pi
 12'b100011111110: begin out_real=16'b1100010011001100; out_imag=16'b1110011110110001; end // in_theta = 1.124023 pi
 12'b100011111111: begin out_real=16'b1100010011010110; out_imag=16'b1110011110011001; end // in_theta = 1.124512 pi
 12'b100100000000: begin out_real=16'b1100010011011111; out_imag=16'b1110011110000010; end // in_theta = 1.125000 pi
 12'b100100000001: begin out_real=16'b1100010011101001; out_imag=16'b1110011101101011; end // in_theta = 1.125488 pi
 12'b100100000010: begin out_real=16'b1100010011110010; out_imag=16'b1110011101010100; end // in_theta = 1.125977 pi
 12'b100100000011: begin out_real=16'b1100010011111100; out_imag=16'b1110011100111101; end // in_theta = 1.126465 pi
 12'b100100000100: begin out_real=16'b1100010100000110; out_imag=16'b1110011100100101; end // in_theta = 1.126953 pi
 12'b100100000101: begin out_real=16'b1100010100010000; out_imag=16'b1110011100001110; end // in_theta = 1.127441 pi
 12'b100100000110: begin out_real=16'b1100010100011010; out_imag=16'b1110011011110111; end // in_theta = 1.127930 pi
 12'b100100000111: begin out_real=16'b1100010100100011; out_imag=16'b1110011011100000; end // in_theta = 1.128418 pi
 12'b100100001000: begin out_real=16'b1100010100101101; out_imag=16'b1110011011001001; end // in_theta = 1.128906 pi
 12'b100100001001: begin out_real=16'b1100010100110111; out_imag=16'b1110011010110010; end // in_theta = 1.129395 pi
 12'b100100001010: begin out_real=16'b1100010101000001; out_imag=16'b1110011010011011; end // in_theta = 1.129883 pi
 12'b100100001011: begin out_real=16'b1100010101001011; out_imag=16'b1110011010000100; end // in_theta = 1.130371 pi
 12'b100100001100: begin out_real=16'b1100010101010101; out_imag=16'b1110011001101101; end // in_theta = 1.130859 pi
 12'b100100001101: begin out_real=16'b1100010101011111; out_imag=16'b1110011001010110; end // in_theta = 1.131348 pi
 12'b100100001110: begin out_real=16'b1100010101101001; out_imag=16'b1110011000111111; end // in_theta = 1.131836 pi
 12'b100100001111: begin out_real=16'b1100010101110011; out_imag=16'b1110011000101000; end // in_theta = 1.132324 pi
 12'b100100010000: begin out_real=16'b1100010101111110; out_imag=16'b1110011000010001; end // in_theta = 1.132813 pi
 12'b100100010001: begin out_real=16'b1100010110001000; out_imag=16'b1110010111111010; end // in_theta = 1.133301 pi
 12'b100100010010: begin out_real=16'b1100010110010010; out_imag=16'b1110010111100011; end // in_theta = 1.133789 pi
 12'b100100010011: begin out_real=16'b1100010110011100; out_imag=16'b1110010111001100; end // in_theta = 1.134277 pi
 12'b100100010100: begin out_real=16'b1100010110100111; out_imag=16'b1110010110110101; end // in_theta = 1.134766 pi
 12'b100100010101: begin out_real=16'b1100010110110001; out_imag=16'b1110010110011110; end // in_theta = 1.135254 pi
 12'b100100010110: begin out_real=16'b1100010110111011; out_imag=16'b1110010110000111; end // in_theta = 1.135742 pi
 12'b100100010111: begin out_real=16'b1100010111000110; out_imag=16'b1110010101110000; end // in_theta = 1.136230 pi
 12'b100100011000: begin out_real=16'b1100010111010000; out_imag=16'b1110010101011001; end // in_theta = 1.136719 pi
 12'b100100011001: begin out_real=16'b1100010111011011; out_imag=16'b1110010101000010; end // in_theta = 1.137207 pi
 12'b100100011010: begin out_real=16'b1100010111100101; out_imag=16'b1110010100101100; end // in_theta = 1.137695 pi
 12'b100100011011: begin out_real=16'b1100010111110000; out_imag=16'b1110010100010101; end // in_theta = 1.138184 pi
 12'b100100011100: begin out_real=16'b1100010111111010; out_imag=16'b1110010011111110; end // in_theta = 1.138672 pi
 12'b100100011101: begin out_real=16'b1100011000000101; out_imag=16'b1110010011100111; end // in_theta = 1.139160 pi
 12'b100100011110: begin out_real=16'b1100011000010000; out_imag=16'b1110010011010000; end // in_theta = 1.139648 pi
 12'b100100011111: begin out_real=16'b1100011000011010; out_imag=16'b1110010010111010; end // in_theta = 1.140137 pi
 12'b100100100000: begin out_real=16'b1100011000100101; out_imag=16'b1110010010100011; end // in_theta = 1.140625 pi
 12'b100100100001: begin out_real=16'b1100011000110000; out_imag=16'b1110010010001100; end // in_theta = 1.141113 pi
 12'b100100100010: begin out_real=16'b1100011000111011; out_imag=16'b1110010001110110; end // in_theta = 1.141602 pi
 12'b100100100011: begin out_real=16'b1100011001000101; out_imag=16'b1110010001011111; end // in_theta = 1.142090 pi
 12'b100100100100: begin out_real=16'b1100011001010000; out_imag=16'b1110010001001000; end // in_theta = 1.142578 pi
 12'b100100100101: begin out_real=16'b1100011001011011; out_imag=16'b1110010000110010; end // in_theta = 1.143066 pi
 12'b100100100110: begin out_real=16'b1100011001100110; out_imag=16'b1110010000011011; end // in_theta = 1.143555 pi
 12'b100100100111: begin out_real=16'b1100011001110001; out_imag=16'b1110010000000100; end // in_theta = 1.144043 pi
 12'b100100101000: begin out_real=16'b1100011001111100; out_imag=16'b1110001111101110; end // in_theta = 1.144531 pi
 12'b100100101001: begin out_real=16'b1100011010000111; out_imag=16'b1110001111010111; end // in_theta = 1.145020 pi
 12'b100100101010: begin out_real=16'b1100011010010010; out_imag=16'b1110001111000001; end // in_theta = 1.145508 pi
 12'b100100101011: begin out_real=16'b1100011010011101; out_imag=16'b1110001110101010; end // in_theta = 1.145996 pi
 12'b100100101100: begin out_real=16'b1100011010101000; out_imag=16'b1110001110010100; end // in_theta = 1.146484 pi
 12'b100100101101: begin out_real=16'b1100011010110100; out_imag=16'b1110001101111101; end // in_theta = 1.146973 pi
 12'b100100101110: begin out_real=16'b1100011010111111; out_imag=16'b1110001101100111; end // in_theta = 1.147461 pi
 12'b100100101111: begin out_real=16'b1100011011001010; out_imag=16'b1110001101010000; end // in_theta = 1.147949 pi
 12'b100100110000: begin out_real=16'b1100011011010101; out_imag=16'b1110001100111010; end // in_theta = 1.148438 pi
 12'b100100110001: begin out_real=16'b1100011011100001; out_imag=16'b1110001100100011; end // in_theta = 1.148926 pi
 12'b100100110010: begin out_real=16'b1100011011101100; out_imag=16'b1110001100001101; end // in_theta = 1.149414 pi
 12'b100100110011: begin out_real=16'b1100011011110111; out_imag=16'b1110001011110110; end // in_theta = 1.149902 pi
 12'b100100110100: begin out_real=16'b1100011100000011; out_imag=16'b1110001011100000; end // in_theta = 1.150391 pi
 12'b100100110101: begin out_real=16'b1100011100001110; out_imag=16'b1110001011001010; end // in_theta = 1.150879 pi
 12'b100100110110: begin out_real=16'b1100011100011010; out_imag=16'b1110001010110011; end // in_theta = 1.151367 pi
 12'b100100110111: begin out_real=16'b1100011100100101; out_imag=16'b1110001010011101; end // in_theta = 1.151855 pi
 12'b100100111000: begin out_real=16'b1100011100110001; out_imag=16'b1110001010000111; end // in_theta = 1.152344 pi
 12'b100100111001: begin out_real=16'b1100011100111101; out_imag=16'b1110001001110000; end // in_theta = 1.152832 pi
 12'b100100111010: begin out_real=16'b1100011101001000; out_imag=16'b1110001001011010; end // in_theta = 1.153320 pi
 12'b100100111011: begin out_real=16'b1100011101010100; out_imag=16'b1110001001000100; end // in_theta = 1.153809 pi
 12'b100100111100: begin out_real=16'b1100011101011111; out_imag=16'b1110001000101101; end // in_theta = 1.154297 pi
 12'b100100111101: begin out_real=16'b1100011101101011; out_imag=16'b1110001000010111; end // in_theta = 1.154785 pi
 12'b100100111110: begin out_real=16'b1100011101110111; out_imag=16'b1110001000000001; end // in_theta = 1.155273 pi
 12'b100100111111: begin out_real=16'b1100011110000011; out_imag=16'b1110000111101011; end // in_theta = 1.155762 pi
 12'b100101000000: begin out_real=16'b1100011110001111; out_imag=16'b1110000111010101; end // in_theta = 1.156250 pi
 12'b100101000001: begin out_real=16'b1100011110011010; out_imag=16'b1110000110111110; end // in_theta = 1.156738 pi
 12'b100101000010: begin out_real=16'b1100011110100110; out_imag=16'b1110000110101000; end // in_theta = 1.157227 pi
 12'b100101000011: begin out_real=16'b1100011110110010; out_imag=16'b1110000110010010; end // in_theta = 1.157715 pi
 12'b100101000100: begin out_real=16'b1100011110111110; out_imag=16'b1110000101111100; end // in_theta = 1.158203 pi
 12'b100101000101: begin out_real=16'b1100011111001010; out_imag=16'b1110000101100110; end // in_theta = 1.158691 pi
 12'b100101000110: begin out_real=16'b1100011111010110; out_imag=16'b1110000101010000; end // in_theta = 1.159180 pi
 12'b100101000111: begin out_real=16'b1100011111100010; out_imag=16'b1110000100111010; end // in_theta = 1.159668 pi
 12'b100101001000: begin out_real=16'b1100011111101110; out_imag=16'b1110000100100100; end // in_theta = 1.160156 pi
 12'b100101001001: begin out_real=16'b1100011111111011; out_imag=16'b1110000100001110; end // in_theta = 1.160645 pi
 12'b100101001010: begin out_real=16'b1100100000000111; out_imag=16'b1110000011111000; end // in_theta = 1.161133 pi
 12'b100101001011: begin out_real=16'b1100100000010011; out_imag=16'b1110000011100010; end // in_theta = 1.161621 pi
 12'b100101001100: begin out_real=16'b1100100000011111; out_imag=16'b1110000011001100; end // in_theta = 1.162109 pi
 12'b100101001101: begin out_real=16'b1100100000101011; out_imag=16'b1110000010110110; end // in_theta = 1.162598 pi
 12'b100101001110: begin out_real=16'b1100100000111000; out_imag=16'b1110000010100000; end // in_theta = 1.163086 pi
 12'b100101001111: begin out_real=16'b1100100001000100; out_imag=16'b1110000010001010; end // in_theta = 1.163574 pi
 12'b100101010000: begin out_real=16'b1100100001010000; out_imag=16'b1110000001110100; end // in_theta = 1.164063 pi
 12'b100101010001: begin out_real=16'b1100100001011101; out_imag=16'b1110000001011110; end // in_theta = 1.164551 pi
 12'b100101010010: begin out_real=16'b1100100001101001; out_imag=16'b1110000001001001; end // in_theta = 1.165039 pi
 12'b100101010011: begin out_real=16'b1100100001110110; out_imag=16'b1110000000110011; end // in_theta = 1.165527 pi
 12'b100101010100: begin out_real=16'b1100100010000010; out_imag=16'b1110000000011101; end // in_theta = 1.166016 pi
 12'b100101010101: begin out_real=16'b1100100010001111; out_imag=16'b1110000000000111; end // in_theta = 1.166504 pi
 12'b100101010110: begin out_real=16'b1100100010011011; out_imag=16'b1101111111110001; end // in_theta = 1.166992 pi
 12'b100101010111: begin out_real=16'b1100100010101000; out_imag=16'b1101111111011100; end // in_theta = 1.167480 pi
 12'b100101011000: begin out_real=16'b1100100010110101; out_imag=16'b1101111111000110; end // in_theta = 1.167969 pi
 12'b100101011001: begin out_real=16'b1100100011000001; out_imag=16'b1101111110110000; end // in_theta = 1.168457 pi
 12'b100101011010: begin out_real=16'b1100100011001110; out_imag=16'b1101111110011011; end // in_theta = 1.168945 pi
 12'b100101011011: begin out_real=16'b1100100011011011; out_imag=16'b1101111110000101; end // in_theta = 1.169434 pi
 12'b100101011100: begin out_real=16'b1100100011101000; out_imag=16'b1101111101101111; end // in_theta = 1.169922 pi
 12'b100101011101: begin out_real=16'b1100100011110100; out_imag=16'b1101111101011010; end // in_theta = 1.170410 pi
 12'b100101011110: begin out_real=16'b1100100100000001; out_imag=16'b1101111101000100; end // in_theta = 1.170898 pi
 12'b100101011111: begin out_real=16'b1100100100001110; out_imag=16'b1101111100101111; end // in_theta = 1.171387 pi
 12'b100101100000: begin out_real=16'b1100100100011011; out_imag=16'b1101111100011001; end // in_theta = 1.171875 pi
 12'b100101100001: begin out_real=16'b1100100100101000; out_imag=16'b1101111100000011; end // in_theta = 1.172363 pi
 12'b100101100010: begin out_real=16'b1100100100110101; out_imag=16'b1101111011101110; end // in_theta = 1.172852 pi
 12'b100101100011: begin out_real=16'b1100100101000010; out_imag=16'b1101111011011000; end // in_theta = 1.173340 pi
 12'b100101100100: begin out_real=16'b1100100101001111; out_imag=16'b1101111011000011; end // in_theta = 1.173828 pi
 12'b100101100101: begin out_real=16'b1100100101011100; out_imag=16'b1101111010101101; end // in_theta = 1.174316 pi
 12'b100101100110: begin out_real=16'b1100100101101001; out_imag=16'b1101111010011000; end // in_theta = 1.174805 pi
 12'b100101100111: begin out_real=16'b1100100101110110; out_imag=16'b1101111010000011; end // in_theta = 1.175293 pi
 12'b100101101000: begin out_real=16'b1100100110000011; out_imag=16'b1101111001101101; end // in_theta = 1.175781 pi
 12'b100101101001: begin out_real=16'b1100100110010001; out_imag=16'b1101111001011000; end // in_theta = 1.176270 pi
 12'b100101101010: begin out_real=16'b1100100110011110; out_imag=16'b1101111001000010; end // in_theta = 1.176758 pi
 12'b100101101011: begin out_real=16'b1100100110101011; out_imag=16'b1101111000101101; end // in_theta = 1.177246 pi
 12'b100101101100: begin out_real=16'b1100100110111000; out_imag=16'b1101111000011000; end // in_theta = 1.177734 pi
 12'b100101101101: begin out_real=16'b1100100111000110; out_imag=16'b1101111000000010; end // in_theta = 1.178223 pi
 12'b100101101110: begin out_real=16'b1100100111010011; out_imag=16'b1101110111101101; end // in_theta = 1.178711 pi
 12'b100101101111: begin out_real=16'b1100100111100000; out_imag=16'b1101110111011000; end // in_theta = 1.179199 pi
 12'b100101110000: begin out_real=16'b1100100111101110; out_imag=16'b1101110111000011; end // in_theta = 1.179688 pi
 12'b100101110001: begin out_real=16'b1100100111111011; out_imag=16'b1101110110101101; end // in_theta = 1.180176 pi
 12'b100101110010: begin out_real=16'b1100101000001001; out_imag=16'b1101110110011000; end // in_theta = 1.180664 pi
 12'b100101110011: begin out_real=16'b1100101000010110; out_imag=16'b1101110110000011; end // in_theta = 1.181152 pi
 12'b100101110100: begin out_real=16'b1100101000100100; out_imag=16'b1101110101101110; end // in_theta = 1.181641 pi
 12'b100101110101: begin out_real=16'b1100101000110010; out_imag=16'b1101110101011001; end // in_theta = 1.182129 pi
 12'b100101110110: begin out_real=16'b1100101000111111; out_imag=16'b1101110101000100; end // in_theta = 1.182617 pi
 12'b100101110111: begin out_real=16'b1100101001001101; out_imag=16'b1101110100101110; end // in_theta = 1.183105 pi
 12'b100101111000: begin out_real=16'b1100101001011011; out_imag=16'b1101110100011001; end // in_theta = 1.183594 pi
 12'b100101111001: begin out_real=16'b1100101001101000; out_imag=16'b1101110100000100; end // in_theta = 1.184082 pi
 12'b100101111010: begin out_real=16'b1100101001110110; out_imag=16'b1101110011101111; end // in_theta = 1.184570 pi
 12'b100101111011: begin out_real=16'b1100101010000100; out_imag=16'b1101110011011010; end // in_theta = 1.185059 pi
 12'b100101111100: begin out_real=16'b1100101010010010; out_imag=16'b1101110011000101; end // in_theta = 1.185547 pi
 12'b100101111101: begin out_real=16'b1100101010011111; out_imag=16'b1101110010110000; end // in_theta = 1.186035 pi
 12'b100101111110: begin out_real=16'b1100101010101101; out_imag=16'b1101110010011011; end // in_theta = 1.186523 pi
 12'b100101111111: begin out_real=16'b1100101010111011; out_imag=16'b1101110010000110; end // in_theta = 1.187012 pi
 12'b100110000000: begin out_real=16'b1100101011001001; out_imag=16'b1101110001110010; end // in_theta = 1.187500 pi
 12'b100110000001: begin out_real=16'b1100101011010111; out_imag=16'b1101110001011101; end // in_theta = 1.187988 pi
 12'b100110000010: begin out_real=16'b1100101011100101; out_imag=16'b1101110001001000; end // in_theta = 1.188477 pi
 12'b100110000011: begin out_real=16'b1100101011110011; out_imag=16'b1101110000110011; end // in_theta = 1.188965 pi
 12'b100110000100: begin out_real=16'b1100101100000001; out_imag=16'b1101110000011110; end // in_theta = 1.189453 pi
 12'b100110000101: begin out_real=16'b1100101100001111; out_imag=16'b1101110000001001; end // in_theta = 1.189941 pi
 12'b100110000110: begin out_real=16'b1100101100011110; out_imag=16'b1101101111110101; end // in_theta = 1.190430 pi
 12'b100110000111: begin out_real=16'b1100101100101100; out_imag=16'b1101101111100000; end // in_theta = 1.190918 pi
 12'b100110001000: begin out_real=16'b1100101100111010; out_imag=16'b1101101111001011; end // in_theta = 1.191406 pi
 12'b100110001001: begin out_real=16'b1100101101001000; out_imag=16'b1101101110110110; end // in_theta = 1.191895 pi
 12'b100110001010: begin out_real=16'b1100101101010110; out_imag=16'b1101101110100010; end // in_theta = 1.192383 pi
 12'b100110001011: begin out_real=16'b1100101101100101; out_imag=16'b1101101110001101; end // in_theta = 1.192871 pi
 12'b100110001100: begin out_real=16'b1100101101110011; out_imag=16'b1101101101111000; end // in_theta = 1.193359 pi
 12'b100110001101: begin out_real=16'b1100101110000001; out_imag=16'b1101101101100100; end // in_theta = 1.193848 pi
 12'b100110001110: begin out_real=16'b1100101110010000; out_imag=16'b1101101101001111; end // in_theta = 1.194336 pi
 12'b100110001111: begin out_real=16'b1100101110011110; out_imag=16'b1101101100111011; end // in_theta = 1.194824 pi
 12'b100110010000: begin out_real=16'b1100101110101101; out_imag=16'b1101101100100110; end // in_theta = 1.195313 pi
 12'b100110010001: begin out_real=16'b1100101110111011; out_imag=16'b1101101100010001; end // in_theta = 1.195801 pi
 12'b100110010010: begin out_real=16'b1100101111001010; out_imag=16'b1101101011111101; end // in_theta = 1.196289 pi
 12'b100110010011: begin out_real=16'b1100101111011000; out_imag=16'b1101101011101000; end // in_theta = 1.196777 pi
 12'b100110010100: begin out_real=16'b1100101111100111; out_imag=16'b1101101011010100; end // in_theta = 1.197266 pi
 12'b100110010101: begin out_real=16'b1100101111110101; out_imag=16'b1101101010111111; end // in_theta = 1.197754 pi
 12'b100110010110: begin out_real=16'b1100110000000100; out_imag=16'b1101101010101011; end // in_theta = 1.198242 pi
 12'b100110010111: begin out_real=16'b1100110000010011; out_imag=16'b1101101010010111; end // in_theta = 1.198730 pi
 12'b100110011000: begin out_real=16'b1100110000100001; out_imag=16'b1101101010000010; end // in_theta = 1.199219 pi
 12'b100110011001: begin out_real=16'b1100110000110000; out_imag=16'b1101101001101110; end // in_theta = 1.199707 pi
 12'b100110011010: begin out_real=16'b1100110000111111; out_imag=16'b1101101001011010; end // in_theta = 1.200195 pi
 12'b100110011011: begin out_real=16'b1100110001001110; out_imag=16'b1101101001000101; end // in_theta = 1.200684 pi
 12'b100110011100: begin out_real=16'b1100110001011101; out_imag=16'b1101101000110001; end // in_theta = 1.201172 pi
 12'b100110011101: begin out_real=16'b1100110001101011; out_imag=16'b1101101000011101; end // in_theta = 1.201660 pi
 12'b100110011110: begin out_real=16'b1100110001111010; out_imag=16'b1101101000001000; end // in_theta = 1.202148 pi
 12'b100110011111: begin out_real=16'b1100110010001001; out_imag=16'b1101100111110100; end // in_theta = 1.202637 pi
 12'b100110100000: begin out_real=16'b1100110010011000; out_imag=16'b1101100111100000; end // in_theta = 1.203125 pi
 12'b100110100001: begin out_real=16'b1100110010100111; out_imag=16'b1101100111001100; end // in_theta = 1.203613 pi
 12'b100110100010: begin out_real=16'b1100110010110110; out_imag=16'b1101100110111000; end // in_theta = 1.204102 pi
 12'b100110100011: begin out_real=16'b1100110011000101; out_imag=16'b1101100110100100; end // in_theta = 1.204590 pi
 12'b100110100100: begin out_real=16'b1100110011010100; out_imag=16'b1101100110001111; end // in_theta = 1.205078 pi
 12'b100110100101: begin out_real=16'b1100110011100011; out_imag=16'b1101100101111011; end // in_theta = 1.205566 pi
 12'b100110100110: begin out_real=16'b1100110011110011; out_imag=16'b1101100101100111; end // in_theta = 1.206055 pi
 12'b100110100111: begin out_real=16'b1100110100000010; out_imag=16'b1101100101010011; end // in_theta = 1.206543 pi
 12'b100110101000: begin out_real=16'b1100110100010001; out_imag=16'b1101100100111111; end // in_theta = 1.207031 pi
 12'b100110101001: begin out_real=16'b1100110100100000; out_imag=16'b1101100100101011; end // in_theta = 1.207520 pi
 12'b100110101010: begin out_real=16'b1100110100110000; out_imag=16'b1101100100010111; end // in_theta = 1.208008 pi
 12'b100110101011: begin out_real=16'b1100110100111111; out_imag=16'b1101100100000011; end // in_theta = 1.208496 pi
 12'b100110101100: begin out_real=16'b1100110101001110; out_imag=16'b1101100011101111; end // in_theta = 1.208984 pi
 12'b100110101101: begin out_real=16'b1100110101011101; out_imag=16'b1101100011011100; end // in_theta = 1.209473 pi
 12'b100110101110: begin out_real=16'b1100110101101101; out_imag=16'b1101100011001000; end // in_theta = 1.209961 pi
 12'b100110101111: begin out_real=16'b1100110101111100; out_imag=16'b1101100010110100; end // in_theta = 1.210449 pi
 12'b100110110000: begin out_real=16'b1100110110001100; out_imag=16'b1101100010100000; end // in_theta = 1.210938 pi
 12'b100110110001: begin out_real=16'b1100110110011011; out_imag=16'b1101100010001100; end // in_theta = 1.211426 pi
 12'b100110110010: begin out_real=16'b1100110110101011; out_imag=16'b1101100001111000; end // in_theta = 1.211914 pi
 12'b100110110011: begin out_real=16'b1100110110111010; out_imag=16'b1101100001100101; end // in_theta = 1.212402 pi
 12'b100110110100: begin out_real=16'b1100110111001010; out_imag=16'b1101100001010001; end // in_theta = 1.212891 pi
 12'b100110110101: begin out_real=16'b1100110111011001; out_imag=16'b1101100000111101; end // in_theta = 1.213379 pi
 12'b100110110110: begin out_real=16'b1100110111101001; out_imag=16'b1101100000101010; end // in_theta = 1.213867 pi
 12'b100110110111: begin out_real=16'b1100110111111001; out_imag=16'b1101100000010110; end // in_theta = 1.214355 pi
 12'b100110111000: begin out_real=16'b1100111000001000; out_imag=16'b1101100000000010; end // in_theta = 1.214844 pi
 12'b100110111001: begin out_real=16'b1100111000011000; out_imag=16'b1101011111101111; end // in_theta = 1.215332 pi
 12'b100110111010: begin out_real=16'b1100111000101000; out_imag=16'b1101011111011011; end // in_theta = 1.215820 pi
 12'b100110111011: begin out_real=16'b1100111000111000; out_imag=16'b1101011111001000; end // in_theta = 1.216309 pi
 12'b100110111100: begin out_real=16'b1100111001000111; out_imag=16'b1101011110110100; end // in_theta = 1.216797 pi
 12'b100110111101: begin out_real=16'b1100111001010111; out_imag=16'b1101011110100000; end // in_theta = 1.217285 pi
 12'b100110111110: begin out_real=16'b1100111001100111; out_imag=16'b1101011110001101; end // in_theta = 1.217773 pi
 12'b100110111111: begin out_real=16'b1100111001110111; out_imag=16'b1101011101111010; end // in_theta = 1.218262 pi
 12'b100111000000: begin out_real=16'b1100111010000111; out_imag=16'b1101011101100110; end // in_theta = 1.218750 pi
 12'b100111000001: begin out_real=16'b1100111010010111; out_imag=16'b1101011101010011; end // in_theta = 1.219238 pi
 12'b100111000010: begin out_real=16'b1100111010100111; out_imag=16'b1101011100111111; end // in_theta = 1.219727 pi
 12'b100111000011: begin out_real=16'b1100111010110111; out_imag=16'b1101011100101100; end // in_theta = 1.220215 pi
 12'b100111000100: begin out_real=16'b1100111011000111; out_imag=16'b1101011100011001; end // in_theta = 1.220703 pi
 12'b100111000101: begin out_real=16'b1100111011010111; out_imag=16'b1101011100000101; end // in_theta = 1.221191 pi
 12'b100111000110: begin out_real=16'b1100111011100111; out_imag=16'b1101011011110010; end // in_theta = 1.221680 pi
 12'b100111000111: begin out_real=16'b1100111011110111; out_imag=16'b1101011011011111; end // in_theta = 1.222168 pi
 12'b100111001000: begin out_real=16'b1100111100000111; out_imag=16'b1101011011001011; end // in_theta = 1.222656 pi
 12'b100111001001: begin out_real=16'b1100111100011000; out_imag=16'b1101011010111000; end // in_theta = 1.223145 pi
 12'b100111001010: begin out_real=16'b1100111100101000; out_imag=16'b1101011010100101; end // in_theta = 1.223633 pi
 12'b100111001011: begin out_real=16'b1100111100111000; out_imag=16'b1101011010010010; end // in_theta = 1.224121 pi
 12'b100111001100: begin out_real=16'b1100111101001000; out_imag=16'b1101011001111111; end // in_theta = 1.224609 pi
 12'b100111001101: begin out_real=16'b1100111101011001; out_imag=16'b1101011001101100; end // in_theta = 1.225098 pi
 12'b100111001110: begin out_real=16'b1100111101101001; out_imag=16'b1101011001011001; end // in_theta = 1.225586 pi
 12'b100111001111: begin out_real=16'b1100111101111001; out_imag=16'b1101011001000101; end // in_theta = 1.226074 pi
 12'b100111010000: begin out_real=16'b1100111110001010; out_imag=16'b1101011000110010; end // in_theta = 1.226563 pi
 12'b100111010001: begin out_real=16'b1100111110011010; out_imag=16'b1101011000011111; end // in_theta = 1.227051 pi
 12'b100111010010: begin out_real=16'b1100111110101011; out_imag=16'b1101011000001100; end // in_theta = 1.227539 pi
 12'b100111010011: begin out_real=16'b1100111110111011; out_imag=16'b1101010111111001; end // in_theta = 1.228027 pi
 12'b100111010100: begin out_real=16'b1100111111001100; out_imag=16'b1101010111100110; end // in_theta = 1.228516 pi
 12'b100111010101: begin out_real=16'b1100111111011100; out_imag=16'b1101010111010100; end // in_theta = 1.229004 pi
 12'b100111010110: begin out_real=16'b1100111111101101; out_imag=16'b1101010111000001; end // in_theta = 1.229492 pi
 12'b100111010111: begin out_real=16'b1100111111111110; out_imag=16'b1101010110101110; end // in_theta = 1.229980 pi
 12'b100111011000: begin out_real=16'b1101000000001110; out_imag=16'b1101010110011011; end // in_theta = 1.230469 pi
 12'b100111011001: begin out_real=16'b1101000000011111; out_imag=16'b1101010110001000; end // in_theta = 1.230957 pi
 12'b100111011010: begin out_real=16'b1101000000110000; out_imag=16'b1101010101110101; end // in_theta = 1.231445 pi
 12'b100111011011: begin out_real=16'b1101000001000000; out_imag=16'b1101010101100011; end // in_theta = 1.231934 pi
 12'b100111011100: begin out_real=16'b1101000001010001; out_imag=16'b1101010101010000; end // in_theta = 1.232422 pi
 12'b100111011101: begin out_real=16'b1101000001100010; out_imag=16'b1101010100111101; end // in_theta = 1.232910 pi
 12'b100111011110: begin out_real=16'b1101000001110011; out_imag=16'b1101010100101010; end // in_theta = 1.233398 pi
 12'b100111011111: begin out_real=16'b1101000010000011; out_imag=16'b1101010100011000; end // in_theta = 1.233887 pi
 12'b100111100000: begin out_real=16'b1101000010010100; out_imag=16'b1101010100000101; end // in_theta = 1.234375 pi
 12'b100111100001: begin out_real=16'b1101000010100101; out_imag=16'b1101010011110011; end // in_theta = 1.234863 pi
 12'b100111100010: begin out_real=16'b1101000010110110; out_imag=16'b1101010011100000; end // in_theta = 1.235352 pi
 12'b100111100011: begin out_real=16'b1101000011000111; out_imag=16'b1101010011001101; end // in_theta = 1.235840 pi
 12'b100111100100: begin out_real=16'b1101000011011000; out_imag=16'b1101010010111011; end // in_theta = 1.236328 pi
 12'b100111100101: begin out_real=16'b1101000011101001; out_imag=16'b1101010010101000; end // in_theta = 1.236816 pi
 12'b100111100110: begin out_real=16'b1101000011111010; out_imag=16'b1101010010010110; end // in_theta = 1.237305 pi
 12'b100111100111: begin out_real=16'b1101000100001011; out_imag=16'b1101010010000011; end // in_theta = 1.237793 pi
 12'b100111101000: begin out_real=16'b1101000100011100; out_imag=16'b1101010001110001; end // in_theta = 1.238281 pi
 12'b100111101001: begin out_real=16'b1101000100101101; out_imag=16'b1101010001011111; end // in_theta = 1.238770 pi
 12'b100111101010: begin out_real=16'b1101000100111110; out_imag=16'b1101010001001100; end // in_theta = 1.239258 pi
 12'b100111101011: begin out_real=16'b1101000101010000; out_imag=16'b1101010000111010; end // in_theta = 1.239746 pi
 12'b100111101100: begin out_real=16'b1101000101100001; out_imag=16'b1101010000101000; end // in_theta = 1.240234 pi
 12'b100111101101: begin out_real=16'b1101000101110010; out_imag=16'b1101010000010101; end // in_theta = 1.240723 pi
 12'b100111101110: begin out_real=16'b1101000110000011; out_imag=16'b1101010000000011; end // in_theta = 1.241211 pi
 12'b100111101111: begin out_real=16'b1101000110010101; out_imag=16'b1101001111110001; end // in_theta = 1.241699 pi
 12'b100111110000: begin out_real=16'b1101000110100110; out_imag=16'b1101001111011111; end // in_theta = 1.242188 pi
 12'b100111110001: begin out_real=16'b1101000110110111; out_imag=16'b1101001111001100; end // in_theta = 1.242676 pi
 12'b100111110010: begin out_real=16'b1101000111001001; out_imag=16'b1101001110111010; end // in_theta = 1.243164 pi
 12'b100111110011: begin out_real=16'b1101000111011010; out_imag=16'b1101001110101000; end // in_theta = 1.243652 pi
 12'b100111110100: begin out_real=16'b1101000111101011; out_imag=16'b1101001110010110; end // in_theta = 1.244141 pi
 12'b100111110101: begin out_real=16'b1101000111111101; out_imag=16'b1101001110000100; end // in_theta = 1.244629 pi
 12'b100111110110: begin out_real=16'b1101001000001110; out_imag=16'b1101001101110010; end // in_theta = 1.245117 pi
 12'b100111110111: begin out_real=16'b1101001000100000; out_imag=16'b1101001101100000; end // in_theta = 1.245605 pi
 12'b100111111000: begin out_real=16'b1101001000110001; out_imag=16'b1101001101001110; end // in_theta = 1.246094 pi
 12'b100111111001: begin out_real=16'b1101001001000011; out_imag=16'b1101001100111100; end // in_theta = 1.246582 pi
 12'b100111111010: begin out_real=16'b1101001001010101; out_imag=16'b1101001100101010; end // in_theta = 1.247070 pi
 12'b100111111011: begin out_real=16'b1101001001100110; out_imag=16'b1101001100011000; end // in_theta = 1.247559 pi
 12'b100111111100: begin out_real=16'b1101001001111000; out_imag=16'b1101001100000110; end // in_theta = 1.248047 pi
 12'b100111111101: begin out_real=16'b1101001010001010; out_imag=16'b1101001011110100; end // in_theta = 1.248535 pi
 12'b100111111110: begin out_real=16'b1101001010011011; out_imag=16'b1101001011100010; end // in_theta = 1.249023 pi
 12'b100111111111: begin out_real=16'b1101001010101101; out_imag=16'b1101001011010001; end // in_theta = 1.249512 pi
 12'b101000000000: begin out_real=16'b1101001010111111; out_imag=16'b1101001010111111; end // in_theta = 1.250000 pi
 12'b101000000001: begin out_real=16'b1101001011010001; out_imag=16'b1101001010101101; end // in_theta = 1.250488 pi
 12'b101000000010: begin out_real=16'b1101001011100010; out_imag=16'b1101001010011011; end // in_theta = 1.250977 pi
 12'b101000000011: begin out_real=16'b1101001011110100; out_imag=16'b1101001010001010; end // in_theta = 1.251465 pi
 12'b101000000100: begin out_real=16'b1101001100000110; out_imag=16'b1101001001111000; end // in_theta = 1.251953 pi
 12'b101000000101: begin out_real=16'b1101001100011000; out_imag=16'b1101001001100110; end // in_theta = 1.252441 pi
 12'b101000000110: begin out_real=16'b1101001100101010; out_imag=16'b1101001001010101; end // in_theta = 1.252930 pi
 12'b101000000111: begin out_real=16'b1101001100111100; out_imag=16'b1101001001000011; end // in_theta = 1.253418 pi
 12'b101000001000: begin out_real=16'b1101001101001110; out_imag=16'b1101001000110001; end // in_theta = 1.253906 pi
 12'b101000001001: begin out_real=16'b1101001101100000; out_imag=16'b1101001000100000; end // in_theta = 1.254395 pi
 12'b101000001010: begin out_real=16'b1101001101110010; out_imag=16'b1101001000001110; end // in_theta = 1.254883 pi
 12'b101000001011: begin out_real=16'b1101001110000100; out_imag=16'b1101000111111101; end // in_theta = 1.255371 pi
 12'b101000001100: begin out_real=16'b1101001110010110; out_imag=16'b1101000111101011; end // in_theta = 1.255859 pi
 12'b101000001101: begin out_real=16'b1101001110101000; out_imag=16'b1101000111011010; end // in_theta = 1.256348 pi
 12'b101000001110: begin out_real=16'b1101001110111010; out_imag=16'b1101000111001001; end // in_theta = 1.256836 pi
 12'b101000001111: begin out_real=16'b1101001111001100; out_imag=16'b1101000110110111; end // in_theta = 1.257324 pi
 12'b101000010000: begin out_real=16'b1101001111011111; out_imag=16'b1101000110100110; end // in_theta = 1.257813 pi
 12'b101000010001: begin out_real=16'b1101001111110001; out_imag=16'b1101000110010101; end // in_theta = 1.258301 pi
 12'b101000010010: begin out_real=16'b1101010000000011; out_imag=16'b1101000110000011; end // in_theta = 1.258789 pi
 12'b101000010011: begin out_real=16'b1101010000010101; out_imag=16'b1101000101110010; end // in_theta = 1.259277 pi
 12'b101000010100: begin out_real=16'b1101010000101000; out_imag=16'b1101000101100001; end // in_theta = 1.259766 pi
 12'b101000010101: begin out_real=16'b1101010000111010; out_imag=16'b1101000101010000; end // in_theta = 1.260254 pi
 12'b101000010110: begin out_real=16'b1101010001001100; out_imag=16'b1101000100111110; end // in_theta = 1.260742 pi
 12'b101000010111: begin out_real=16'b1101010001011111; out_imag=16'b1101000100101101; end // in_theta = 1.261230 pi
 12'b101000011000: begin out_real=16'b1101010001110001; out_imag=16'b1101000100011100; end // in_theta = 1.261719 pi
 12'b101000011001: begin out_real=16'b1101010010000011; out_imag=16'b1101000100001011; end // in_theta = 1.262207 pi
 12'b101000011010: begin out_real=16'b1101010010010110; out_imag=16'b1101000011111010; end // in_theta = 1.262695 pi
 12'b101000011011: begin out_real=16'b1101010010101000; out_imag=16'b1101000011101001; end // in_theta = 1.263184 pi
 12'b101000011100: begin out_real=16'b1101010010111011; out_imag=16'b1101000011011000; end // in_theta = 1.263672 pi
 12'b101000011101: begin out_real=16'b1101010011001101; out_imag=16'b1101000011000111; end // in_theta = 1.264160 pi
 12'b101000011110: begin out_real=16'b1101010011100000; out_imag=16'b1101000010110110; end // in_theta = 1.264648 pi
 12'b101000011111: begin out_real=16'b1101010011110011; out_imag=16'b1101000010100101; end // in_theta = 1.265137 pi
 12'b101000100000: begin out_real=16'b1101010100000101; out_imag=16'b1101000010010100; end // in_theta = 1.265625 pi
 12'b101000100001: begin out_real=16'b1101010100011000; out_imag=16'b1101000010000011; end // in_theta = 1.266113 pi
 12'b101000100010: begin out_real=16'b1101010100101010; out_imag=16'b1101000001110011; end // in_theta = 1.266602 pi
 12'b101000100011: begin out_real=16'b1101010100111101; out_imag=16'b1101000001100010; end // in_theta = 1.267090 pi
 12'b101000100100: begin out_real=16'b1101010101010000; out_imag=16'b1101000001010001; end // in_theta = 1.267578 pi
 12'b101000100101: begin out_real=16'b1101010101100011; out_imag=16'b1101000001000000; end // in_theta = 1.268066 pi
 12'b101000100110: begin out_real=16'b1101010101110101; out_imag=16'b1101000000110000; end // in_theta = 1.268555 pi
 12'b101000100111: begin out_real=16'b1101010110001000; out_imag=16'b1101000000011111; end // in_theta = 1.269043 pi
 12'b101000101000: begin out_real=16'b1101010110011011; out_imag=16'b1101000000001110; end // in_theta = 1.269531 pi
 12'b101000101001: begin out_real=16'b1101010110101110; out_imag=16'b1100111111111110; end // in_theta = 1.270020 pi
 12'b101000101010: begin out_real=16'b1101010111000001; out_imag=16'b1100111111101101; end // in_theta = 1.270508 pi
 12'b101000101011: begin out_real=16'b1101010111010100; out_imag=16'b1100111111011100; end // in_theta = 1.270996 pi
 12'b101000101100: begin out_real=16'b1101010111100110; out_imag=16'b1100111111001100; end // in_theta = 1.271484 pi
 12'b101000101101: begin out_real=16'b1101010111111001; out_imag=16'b1100111110111011; end // in_theta = 1.271973 pi
 12'b101000101110: begin out_real=16'b1101011000001100; out_imag=16'b1100111110101011; end // in_theta = 1.272461 pi
 12'b101000101111: begin out_real=16'b1101011000011111; out_imag=16'b1100111110011010; end // in_theta = 1.272949 pi
 12'b101000110000: begin out_real=16'b1101011000110010; out_imag=16'b1100111110001010; end // in_theta = 1.273438 pi
 12'b101000110001: begin out_real=16'b1101011001000101; out_imag=16'b1100111101111001; end // in_theta = 1.273926 pi
 12'b101000110010: begin out_real=16'b1101011001011001; out_imag=16'b1100111101101001; end // in_theta = 1.274414 pi
 12'b101000110011: begin out_real=16'b1101011001101100; out_imag=16'b1100111101011001; end // in_theta = 1.274902 pi
 12'b101000110100: begin out_real=16'b1101011001111111; out_imag=16'b1100111101001000; end // in_theta = 1.275391 pi
 12'b101000110101: begin out_real=16'b1101011010010010; out_imag=16'b1100111100111000; end // in_theta = 1.275879 pi
 12'b101000110110: begin out_real=16'b1101011010100101; out_imag=16'b1100111100101000; end // in_theta = 1.276367 pi
 12'b101000110111: begin out_real=16'b1101011010111000; out_imag=16'b1100111100011000; end // in_theta = 1.276855 pi
 12'b101000111000: begin out_real=16'b1101011011001011; out_imag=16'b1100111100000111; end // in_theta = 1.277344 pi
 12'b101000111001: begin out_real=16'b1101011011011111; out_imag=16'b1100111011110111; end // in_theta = 1.277832 pi
 12'b101000111010: begin out_real=16'b1101011011110010; out_imag=16'b1100111011100111; end // in_theta = 1.278320 pi
 12'b101000111011: begin out_real=16'b1101011100000101; out_imag=16'b1100111011010111; end // in_theta = 1.278809 pi
 12'b101000111100: begin out_real=16'b1101011100011001; out_imag=16'b1100111011000111; end // in_theta = 1.279297 pi
 12'b101000111101: begin out_real=16'b1101011100101100; out_imag=16'b1100111010110111; end // in_theta = 1.279785 pi
 12'b101000111110: begin out_real=16'b1101011100111111; out_imag=16'b1100111010100111; end // in_theta = 1.280273 pi
 12'b101000111111: begin out_real=16'b1101011101010011; out_imag=16'b1100111010010111; end // in_theta = 1.280762 pi
 12'b101001000000: begin out_real=16'b1101011101100110; out_imag=16'b1100111010000111; end // in_theta = 1.281250 pi
 12'b101001000001: begin out_real=16'b1101011101111010; out_imag=16'b1100111001110111; end // in_theta = 1.281738 pi
 12'b101001000010: begin out_real=16'b1101011110001101; out_imag=16'b1100111001100111; end // in_theta = 1.282227 pi
 12'b101001000011: begin out_real=16'b1101011110100000; out_imag=16'b1100111001010111; end // in_theta = 1.282715 pi
 12'b101001000100: begin out_real=16'b1101011110110100; out_imag=16'b1100111001000111; end // in_theta = 1.283203 pi
 12'b101001000101: begin out_real=16'b1101011111001000; out_imag=16'b1100111000111000; end // in_theta = 1.283691 pi
 12'b101001000110: begin out_real=16'b1101011111011011; out_imag=16'b1100111000101000; end // in_theta = 1.284180 pi
 12'b101001000111: begin out_real=16'b1101011111101111; out_imag=16'b1100111000011000; end // in_theta = 1.284668 pi
 12'b101001001000: begin out_real=16'b1101100000000010; out_imag=16'b1100111000001000; end // in_theta = 1.285156 pi
 12'b101001001001: begin out_real=16'b1101100000010110; out_imag=16'b1100110111111001; end // in_theta = 1.285645 pi
 12'b101001001010: begin out_real=16'b1101100000101010; out_imag=16'b1100110111101001; end // in_theta = 1.286133 pi
 12'b101001001011: begin out_real=16'b1101100000111101; out_imag=16'b1100110111011001; end // in_theta = 1.286621 pi
 12'b101001001100: begin out_real=16'b1101100001010001; out_imag=16'b1100110111001010; end // in_theta = 1.287109 pi
 12'b101001001101: begin out_real=16'b1101100001100101; out_imag=16'b1100110110111010; end // in_theta = 1.287598 pi
 12'b101001001110: begin out_real=16'b1101100001111000; out_imag=16'b1100110110101011; end // in_theta = 1.288086 pi
 12'b101001001111: begin out_real=16'b1101100010001100; out_imag=16'b1100110110011011; end // in_theta = 1.288574 pi
 12'b101001010000: begin out_real=16'b1101100010100000; out_imag=16'b1100110110001100; end // in_theta = 1.289062 pi
 12'b101001010001: begin out_real=16'b1101100010110100; out_imag=16'b1100110101111100; end // in_theta = 1.289551 pi
 12'b101001010010: begin out_real=16'b1101100011001000; out_imag=16'b1100110101101101; end // in_theta = 1.290039 pi
 12'b101001010011: begin out_real=16'b1101100011011100; out_imag=16'b1100110101011101; end // in_theta = 1.290527 pi
 12'b101001010100: begin out_real=16'b1101100011101111; out_imag=16'b1100110101001110; end // in_theta = 1.291016 pi
 12'b101001010101: begin out_real=16'b1101100100000011; out_imag=16'b1100110100111111; end // in_theta = 1.291504 pi
 12'b101001010110: begin out_real=16'b1101100100010111; out_imag=16'b1100110100110000; end // in_theta = 1.291992 pi
 12'b101001010111: begin out_real=16'b1101100100101011; out_imag=16'b1100110100100000; end // in_theta = 1.292480 pi
 12'b101001011000: begin out_real=16'b1101100100111111; out_imag=16'b1100110100010001; end // in_theta = 1.292969 pi
 12'b101001011001: begin out_real=16'b1101100101010011; out_imag=16'b1100110100000010; end // in_theta = 1.293457 pi
 12'b101001011010: begin out_real=16'b1101100101100111; out_imag=16'b1100110011110011; end // in_theta = 1.293945 pi
 12'b101001011011: begin out_real=16'b1101100101111011; out_imag=16'b1100110011100011; end // in_theta = 1.294434 pi
 12'b101001011100: begin out_real=16'b1101100110001111; out_imag=16'b1100110011010100; end // in_theta = 1.294922 pi
 12'b101001011101: begin out_real=16'b1101100110100100; out_imag=16'b1100110011000101; end // in_theta = 1.295410 pi
 12'b101001011110: begin out_real=16'b1101100110111000; out_imag=16'b1100110010110110; end // in_theta = 1.295898 pi
 12'b101001011111: begin out_real=16'b1101100111001100; out_imag=16'b1100110010100111; end // in_theta = 1.296387 pi
 12'b101001100000: begin out_real=16'b1101100111100000; out_imag=16'b1100110010011000; end // in_theta = 1.296875 pi
 12'b101001100001: begin out_real=16'b1101100111110100; out_imag=16'b1100110010001001; end // in_theta = 1.297363 pi
 12'b101001100010: begin out_real=16'b1101101000001000; out_imag=16'b1100110001111010; end // in_theta = 1.297852 pi
 12'b101001100011: begin out_real=16'b1101101000011101; out_imag=16'b1100110001101011; end // in_theta = 1.298340 pi
 12'b101001100100: begin out_real=16'b1101101000110001; out_imag=16'b1100110001011101; end // in_theta = 1.298828 pi
 12'b101001100101: begin out_real=16'b1101101001000101; out_imag=16'b1100110001001110; end // in_theta = 1.299316 pi
 12'b101001100110: begin out_real=16'b1101101001011010; out_imag=16'b1100110000111111; end // in_theta = 1.299805 pi
 12'b101001100111: begin out_real=16'b1101101001101110; out_imag=16'b1100110000110000; end // in_theta = 1.300293 pi
 12'b101001101000: begin out_real=16'b1101101010000010; out_imag=16'b1100110000100001; end // in_theta = 1.300781 pi
 12'b101001101001: begin out_real=16'b1101101010010111; out_imag=16'b1100110000010011; end // in_theta = 1.301270 pi
 12'b101001101010: begin out_real=16'b1101101010101011; out_imag=16'b1100110000000100; end // in_theta = 1.301758 pi
 12'b101001101011: begin out_real=16'b1101101010111111; out_imag=16'b1100101111110101; end // in_theta = 1.302246 pi
 12'b101001101100: begin out_real=16'b1101101011010100; out_imag=16'b1100101111100111; end // in_theta = 1.302734 pi
 12'b101001101101: begin out_real=16'b1101101011101000; out_imag=16'b1100101111011000; end // in_theta = 1.303223 pi
 12'b101001101110: begin out_real=16'b1101101011111101; out_imag=16'b1100101111001010; end // in_theta = 1.303711 pi
 12'b101001101111: begin out_real=16'b1101101100010001; out_imag=16'b1100101110111011; end // in_theta = 1.304199 pi
 12'b101001110000: begin out_real=16'b1101101100100110; out_imag=16'b1100101110101101; end // in_theta = 1.304688 pi
 12'b101001110001: begin out_real=16'b1101101100111011; out_imag=16'b1100101110011110; end // in_theta = 1.305176 pi
 12'b101001110010: begin out_real=16'b1101101101001111; out_imag=16'b1100101110010000; end // in_theta = 1.305664 pi
 12'b101001110011: begin out_real=16'b1101101101100100; out_imag=16'b1100101110000001; end // in_theta = 1.306152 pi
 12'b101001110100: begin out_real=16'b1101101101111000; out_imag=16'b1100101101110011; end // in_theta = 1.306641 pi
 12'b101001110101: begin out_real=16'b1101101110001101; out_imag=16'b1100101101100101; end // in_theta = 1.307129 pi
 12'b101001110110: begin out_real=16'b1101101110100010; out_imag=16'b1100101101010110; end // in_theta = 1.307617 pi
 12'b101001110111: begin out_real=16'b1101101110110110; out_imag=16'b1100101101001000; end // in_theta = 1.308105 pi
 12'b101001111000: begin out_real=16'b1101101111001011; out_imag=16'b1100101100111010; end // in_theta = 1.308594 pi
 12'b101001111001: begin out_real=16'b1101101111100000; out_imag=16'b1100101100101100; end // in_theta = 1.309082 pi
 12'b101001111010: begin out_real=16'b1101101111110101; out_imag=16'b1100101100011110; end // in_theta = 1.309570 pi
 12'b101001111011: begin out_real=16'b1101110000001001; out_imag=16'b1100101100001111; end // in_theta = 1.310059 pi
 12'b101001111100: begin out_real=16'b1101110000011110; out_imag=16'b1100101100000001; end // in_theta = 1.310547 pi
 12'b101001111101: begin out_real=16'b1101110000110011; out_imag=16'b1100101011110011; end // in_theta = 1.311035 pi
 12'b101001111110: begin out_real=16'b1101110001001000; out_imag=16'b1100101011100101; end // in_theta = 1.311523 pi
 12'b101001111111: begin out_real=16'b1101110001011101; out_imag=16'b1100101011010111; end // in_theta = 1.312012 pi
 12'b101010000000: begin out_real=16'b1101110001110010; out_imag=16'b1100101011001001; end // in_theta = 1.312500 pi
 12'b101010000001: begin out_real=16'b1101110010000110; out_imag=16'b1100101010111011; end // in_theta = 1.312988 pi
 12'b101010000010: begin out_real=16'b1101110010011011; out_imag=16'b1100101010101101; end // in_theta = 1.313477 pi
 12'b101010000011: begin out_real=16'b1101110010110000; out_imag=16'b1100101010011111; end // in_theta = 1.313965 pi
 12'b101010000100: begin out_real=16'b1101110011000101; out_imag=16'b1100101010010010; end // in_theta = 1.314453 pi
 12'b101010000101: begin out_real=16'b1101110011011010; out_imag=16'b1100101010000100; end // in_theta = 1.314941 pi
 12'b101010000110: begin out_real=16'b1101110011101111; out_imag=16'b1100101001110110; end // in_theta = 1.315430 pi
 12'b101010000111: begin out_real=16'b1101110100000100; out_imag=16'b1100101001101000; end // in_theta = 1.315918 pi
 12'b101010001000: begin out_real=16'b1101110100011001; out_imag=16'b1100101001011011; end // in_theta = 1.316406 pi
 12'b101010001001: begin out_real=16'b1101110100101110; out_imag=16'b1100101001001101; end // in_theta = 1.316895 pi
 12'b101010001010: begin out_real=16'b1101110101000100; out_imag=16'b1100101000111111; end // in_theta = 1.317383 pi
 12'b101010001011: begin out_real=16'b1101110101011001; out_imag=16'b1100101000110010; end // in_theta = 1.317871 pi
 12'b101010001100: begin out_real=16'b1101110101101110; out_imag=16'b1100101000100100; end // in_theta = 1.318359 pi
 12'b101010001101: begin out_real=16'b1101110110000011; out_imag=16'b1100101000010110; end // in_theta = 1.318848 pi
 12'b101010001110: begin out_real=16'b1101110110011000; out_imag=16'b1100101000001001; end // in_theta = 1.319336 pi
 12'b101010001111: begin out_real=16'b1101110110101101; out_imag=16'b1100100111111011; end // in_theta = 1.319824 pi
 12'b101010010000: begin out_real=16'b1101110111000011; out_imag=16'b1100100111101110; end // in_theta = 1.320313 pi
 12'b101010010001: begin out_real=16'b1101110111011000; out_imag=16'b1100100111100000; end // in_theta = 1.320801 pi
 12'b101010010010: begin out_real=16'b1101110111101101; out_imag=16'b1100100111010011; end // in_theta = 1.321289 pi
 12'b101010010011: begin out_real=16'b1101111000000010; out_imag=16'b1100100111000110; end // in_theta = 1.321777 pi
 12'b101010010100: begin out_real=16'b1101111000011000; out_imag=16'b1100100110111000; end // in_theta = 1.322266 pi
 12'b101010010101: begin out_real=16'b1101111000101101; out_imag=16'b1100100110101011; end // in_theta = 1.322754 pi
 12'b101010010110: begin out_real=16'b1101111001000010; out_imag=16'b1100100110011110; end // in_theta = 1.323242 pi
 12'b101010010111: begin out_real=16'b1101111001011000; out_imag=16'b1100100110010001; end // in_theta = 1.323730 pi
 12'b101010011000: begin out_real=16'b1101111001101101; out_imag=16'b1100100110000011; end // in_theta = 1.324219 pi
 12'b101010011001: begin out_real=16'b1101111010000011; out_imag=16'b1100100101110110; end // in_theta = 1.324707 pi
 12'b101010011010: begin out_real=16'b1101111010011000; out_imag=16'b1100100101101001; end // in_theta = 1.325195 pi
 12'b101010011011: begin out_real=16'b1101111010101101; out_imag=16'b1100100101011100; end // in_theta = 1.325684 pi
 12'b101010011100: begin out_real=16'b1101111011000011; out_imag=16'b1100100101001111; end // in_theta = 1.326172 pi
 12'b101010011101: begin out_real=16'b1101111011011000; out_imag=16'b1100100101000010; end // in_theta = 1.326660 pi
 12'b101010011110: begin out_real=16'b1101111011101110; out_imag=16'b1100100100110101; end // in_theta = 1.327148 pi
 12'b101010011111: begin out_real=16'b1101111100000011; out_imag=16'b1100100100101000; end // in_theta = 1.327637 pi
 12'b101010100000: begin out_real=16'b1101111100011001; out_imag=16'b1100100100011011; end // in_theta = 1.328125 pi
 12'b101010100001: begin out_real=16'b1101111100101111; out_imag=16'b1100100100001110; end // in_theta = 1.328613 pi
 12'b101010100010: begin out_real=16'b1101111101000100; out_imag=16'b1100100100000001; end // in_theta = 1.329102 pi
 12'b101010100011: begin out_real=16'b1101111101011010; out_imag=16'b1100100011110100; end // in_theta = 1.329590 pi
 12'b101010100100: begin out_real=16'b1101111101101111; out_imag=16'b1100100011101000; end // in_theta = 1.330078 pi
 12'b101010100101: begin out_real=16'b1101111110000101; out_imag=16'b1100100011011011; end // in_theta = 1.330566 pi
 12'b101010100110: begin out_real=16'b1101111110011011; out_imag=16'b1100100011001110; end // in_theta = 1.331055 pi
 12'b101010100111: begin out_real=16'b1101111110110000; out_imag=16'b1100100011000001; end // in_theta = 1.331543 pi
 12'b101010101000: begin out_real=16'b1101111111000110; out_imag=16'b1100100010110101; end // in_theta = 1.332031 pi
 12'b101010101001: begin out_real=16'b1101111111011100; out_imag=16'b1100100010101000; end // in_theta = 1.332520 pi
 12'b101010101010: begin out_real=16'b1101111111110001; out_imag=16'b1100100010011011; end // in_theta = 1.333008 pi
 12'b101010101011: begin out_real=16'b1110000000000111; out_imag=16'b1100100010001111; end // in_theta = 1.333496 pi
 12'b101010101100: begin out_real=16'b1110000000011101; out_imag=16'b1100100010000010; end // in_theta = 1.333984 pi
 12'b101010101101: begin out_real=16'b1110000000110011; out_imag=16'b1100100001110110; end // in_theta = 1.334473 pi
 12'b101010101110: begin out_real=16'b1110000001001001; out_imag=16'b1100100001101001; end // in_theta = 1.334961 pi
 12'b101010101111: begin out_real=16'b1110000001011110; out_imag=16'b1100100001011101; end // in_theta = 1.335449 pi
 12'b101010110000: begin out_real=16'b1110000001110100; out_imag=16'b1100100001010000; end // in_theta = 1.335938 pi
 12'b101010110001: begin out_real=16'b1110000010001010; out_imag=16'b1100100001000100; end // in_theta = 1.336426 pi
 12'b101010110010: begin out_real=16'b1110000010100000; out_imag=16'b1100100000111000; end // in_theta = 1.336914 pi
 12'b101010110011: begin out_real=16'b1110000010110110; out_imag=16'b1100100000101011; end // in_theta = 1.337402 pi
 12'b101010110100: begin out_real=16'b1110000011001100; out_imag=16'b1100100000011111; end // in_theta = 1.337891 pi
 12'b101010110101: begin out_real=16'b1110000011100010; out_imag=16'b1100100000010011; end // in_theta = 1.338379 pi
 12'b101010110110: begin out_real=16'b1110000011111000; out_imag=16'b1100100000000111; end // in_theta = 1.338867 pi
 12'b101010110111: begin out_real=16'b1110000100001110; out_imag=16'b1100011111111011; end // in_theta = 1.339355 pi
 12'b101010111000: begin out_real=16'b1110000100100100; out_imag=16'b1100011111101110; end // in_theta = 1.339844 pi
 12'b101010111001: begin out_real=16'b1110000100111010; out_imag=16'b1100011111100010; end // in_theta = 1.340332 pi
 12'b101010111010: begin out_real=16'b1110000101010000; out_imag=16'b1100011111010110; end // in_theta = 1.340820 pi
 12'b101010111011: begin out_real=16'b1110000101100110; out_imag=16'b1100011111001010; end // in_theta = 1.341309 pi
 12'b101010111100: begin out_real=16'b1110000101111100; out_imag=16'b1100011110111110; end // in_theta = 1.341797 pi
 12'b101010111101: begin out_real=16'b1110000110010010; out_imag=16'b1100011110110010; end // in_theta = 1.342285 pi
 12'b101010111110: begin out_real=16'b1110000110101000; out_imag=16'b1100011110100110; end // in_theta = 1.342773 pi
 12'b101010111111: begin out_real=16'b1110000110111110; out_imag=16'b1100011110011010; end // in_theta = 1.343262 pi
 12'b101011000000: begin out_real=16'b1110000111010101; out_imag=16'b1100011110001111; end // in_theta = 1.343750 pi
 12'b101011000001: begin out_real=16'b1110000111101011; out_imag=16'b1100011110000011; end // in_theta = 1.344238 pi
 12'b101011000010: begin out_real=16'b1110001000000001; out_imag=16'b1100011101110111; end // in_theta = 1.344727 pi
 12'b101011000011: begin out_real=16'b1110001000010111; out_imag=16'b1100011101101011; end // in_theta = 1.345215 pi
 12'b101011000100: begin out_real=16'b1110001000101101; out_imag=16'b1100011101011111; end // in_theta = 1.345703 pi
 12'b101011000101: begin out_real=16'b1110001001000100; out_imag=16'b1100011101010100; end // in_theta = 1.346191 pi
 12'b101011000110: begin out_real=16'b1110001001011010; out_imag=16'b1100011101001000; end // in_theta = 1.346680 pi
 12'b101011000111: begin out_real=16'b1110001001110000; out_imag=16'b1100011100111101; end // in_theta = 1.347168 pi
 12'b101011001000: begin out_real=16'b1110001010000111; out_imag=16'b1100011100110001; end // in_theta = 1.347656 pi
 12'b101011001001: begin out_real=16'b1110001010011101; out_imag=16'b1100011100100101; end // in_theta = 1.348145 pi
 12'b101011001010: begin out_real=16'b1110001010110011; out_imag=16'b1100011100011010; end // in_theta = 1.348633 pi
 12'b101011001011: begin out_real=16'b1110001011001010; out_imag=16'b1100011100001110; end // in_theta = 1.349121 pi
 12'b101011001100: begin out_real=16'b1110001011100000; out_imag=16'b1100011100000011; end // in_theta = 1.349609 pi
 12'b101011001101: begin out_real=16'b1110001011110110; out_imag=16'b1100011011110111; end // in_theta = 1.350098 pi
 12'b101011001110: begin out_real=16'b1110001100001101; out_imag=16'b1100011011101100; end // in_theta = 1.350586 pi
 12'b101011001111: begin out_real=16'b1110001100100011; out_imag=16'b1100011011100001; end // in_theta = 1.351074 pi
 12'b101011010000: begin out_real=16'b1110001100111010; out_imag=16'b1100011011010101; end // in_theta = 1.351563 pi
 12'b101011010001: begin out_real=16'b1110001101010000; out_imag=16'b1100011011001010; end // in_theta = 1.352051 pi
 12'b101011010010: begin out_real=16'b1110001101100111; out_imag=16'b1100011010111111; end // in_theta = 1.352539 pi
 12'b101011010011: begin out_real=16'b1110001101111101; out_imag=16'b1100011010110100; end // in_theta = 1.353027 pi
 12'b101011010100: begin out_real=16'b1110001110010100; out_imag=16'b1100011010101000; end // in_theta = 1.353516 pi
 12'b101011010101: begin out_real=16'b1110001110101010; out_imag=16'b1100011010011101; end // in_theta = 1.354004 pi
 12'b101011010110: begin out_real=16'b1110001111000001; out_imag=16'b1100011010010010; end // in_theta = 1.354492 pi
 12'b101011010111: begin out_real=16'b1110001111010111; out_imag=16'b1100011010000111; end // in_theta = 1.354980 pi
 12'b101011011000: begin out_real=16'b1110001111101110; out_imag=16'b1100011001111100; end // in_theta = 1.355469 pi
 12'b101011011001: begin out_real=16'b1110010000000100; out_imag=16'b1100011001110001; end // in_theta = 1.355957 pi
 12'b101011011010: begin out_real=16'b1110010000011011; out_imag=16'b1100011001100110; end // in_theta = 1.356445 pi
 12'b101011011011: begin out_real=16'b1110010000110010; out_imag=16'b1100011001011011; end // in_theta = 1.356934 pi
 12'b101011011100: begin out_real=16'b1110010001001000; out_imag=16'b1100011001010000; end // in_theta = 1.357422 pi
 12'b101011011101: begin out_real=16'b1110010001011111; out_imag=16'b1100011001000101; end // in_theta = 1.357910 pi
 12'b101011011110: begin out_real=16'b1110010001110110; out_imag=16'b1100011000111011; end // in_theta = 1.358398 pi
 12'b101011011111: begin out_real=16'b1110010010001100; out_imag=16'b1100011000110000; end // in_theta = 1.358887 pi
 12'b101011100000: begin out_real=16'b1110010010100011; out_imag=16'b1100011000100101; end // in_theta = 1.359375 pi
 12'b101011100001: begin out_real=16'b1110010010111010; out_imag=16'b1100011000011010; end // in_theta = 1.359863 pi
 12'b101011100010: begin out_real=16'b1110010011010000; out_imag=16'b1100011000010000; end // in_theta = 1.360352 pi
 12'b101011100011: begin out_real=16'b1110010011100111; out_imag=16'b1100011000000101; end // in_theta = 1.360840 pi
 12'b101011100100: begin out_real=16'b1110010011111110; out_imag=16'b1100010111111010; end // in_theta = 1.361328 pi
 12'b101011100101: begin out_real=16'b1110010100010101; out_imag=16'b1100010111110000; end // in_theta = 1.361816 pi
 12'b101011100110: begin out_real=16'b1110010100101100; out_imag=16'b1100010111100101; end // in_theta = 1.362305 pi
 12'b101011100111: begin out_real=16'b1110010101000010; out_imag=16'b1100010111011011; end // in_theta = 1.362793 pi
 12'b101011101000: begin out_real=16'b1110010101011001; out_imag=16'b1100010111010000; end // in_theta = 1.363281 pi
 12'b101011101001: begin out_real=16'b1110010101110000; out_imag=16'b1100010111000110; end // in_theta = 1.363770 pi
 12'b101011101010: begin out_real=16'b1110010110000111; out_imag=16'b1100010110111011; end // in_theta = 1.364258 pi
 12'b101011101011: begin out_real=16'b1110010110011110; out_imag=16'b1100010110110001; end // in_theta = 1.364746 pi
 12'b101011101100: begin out_real=16'b1110010110110101; out_imag=16'b1100010110100111; end // in_theta = 1.365234 pi
 12'b101011101101: begin out_real=16'b1110010111001100; out_imag=16'b1100010110011100; end // in_theta = 1.365723 pi
 12'b101011101110: begin out_real=16'b1110010111100011; out_imag=16'b1100010110010010; end // in_theta = 1.366211 pi
 12'b101011101111: begin out_real=16'b1110010111111010; out_imag=16'b1100010110001000; end // in_theta = 1.366699 pi
 12'b101011110000: begin out_real=16'b1110011000010001; out_imag=16'b1100010101111110; end // in_theta = 1.367187 pi
 12'b101011110001: begin out_real=16'b1110011000101000; out_imag=16'b1100010101110011; end // in_theta = 1.367676 pi
 12'b101011110010: begin out_real=16'b1110011000111111; out_imag=16'b1100010101101001; end // in_theta = 1.368164 pi
 12'b101011110011: begin out_real=16'b1110011001010110; out_imag=16'b1100010101011111; end // in_theta = 1.368652 pi
 12'b101011110100: begin out_real=16'b1110011001101101; out_imag=16'b1100010101010101; end // in_theta = 1.369141 pi
 12'b101011110101: begin out_real=16'b1110011010000100; out_imag=16'b1100010101001011; end // in_theta = 1.369629 pi
 12'b101011110110: begin out_real=16'b1110011010011011; out_imag=16'b1100010101000001; end // in_theta = 1.370117 pi
 12'b101011110111: begin out_real=16'b1110011010110010; out_imag=16'b1100010100110111; end // in_theta = 1.370605 pi
 12'b101011111000: begin out_real=16'b1110011011001001; out_imag=16'b1100010100101101; end // in_theta = 1.371094 pi
 12'b101011111001: begin out_real=16'b1110011011100000; out_imag=16'b1100010100100011; end // in_theta = 1.371582 pi
 12'b101011111010: begin out_real=16'b1110011011110111; out_imag=16'b1100010100011010; end // in_theta = 1.372070 pi
 12'b101011111011: begin out_real=16'b1110011100001110; out_imag=16'b1100010100010000; end // in_theta = 1.372559 pi
 12'b101011111100: begin out_real=16'b1110011100100101; out_imag=16'b1100010100000110; end // in_theta = 1.373047 pi
 12'b101011111101: begin out_real=16'b1110011100111101; out_imag=16'b1100010011111100; end // in_theta = 1.373535 pi
 12'b101011111110: begin out_real=16'b1110011101010100; out_imag=16'b1100010011110010; end // in_theta = 1.374023 pi
 12'b101011111111: begin out_real=16'b1110011101101011; out_imag=16'b1100010011101001; end // in_theta = 1.374512 pi
 12'b101100000000: begin out_real=16'b1110011110000010; out_imag=16'b1100010011011111; end // in_theta = 1.375000 pi
 12'b101100000001: begin out_real=16'b1110011110011001; out_imag=16'b1100010011010110; end // in_theta = 1.375488 pi
 12'b101100000010: begin out_real=16'b1110011110110001; out_imag=16'b1100010011001100; end // in_theta = 1.375977 pi
 12'b101100000011: begin out_real=16'b1110011111001000; out_imag=16'b1100010011000010; end // in_theta = 1.376465 pi
 12'b101100000100: begin out_real=16'b1110011111011111; out_imag=16'b1100010010111001; end // in_theta = 1.376953 pi
 12'b101100000101: begin out_real=16'b1110011111110110; out_imag=16'b1100010010110000; end // in_theta = 1.377441 pi
 12'b101100000110: begin out_real=16'b1110100000001110; out_imag=16'b1100010010100110; end // in_theta = 1.377930 pi
 12'b101100000111: begin out_real=16'b1110100000100101; out_imag=16'b1100010010011101; end // in_theta = 1.378418 pi
 12'b101100001000: begin out_real=16'b1110100000111100; out_imag=16'b1100010010010011; end // in_theta = 1.378906 pi
 12'b101100001001: begin out_real=16'b1110100001010100; out_imag=16'b1100010010001010; end // in_theta = 1.379395 pi
 12'b101100001010: begin out_real=16'b1110100001101011; out_imag=16'b1100010010000001; end // in_theta = 1.379883 pi
 12'b101100001011: begin out_real=16'b1110100010000010; out_imag=16'b1100010001111000; end // in_theta = 1.380371 pi
 12'b101100001100: begin out_real=16'b1110100010011010; out_imag=16'b1100010001101110; end // in_theta = 1.380859 pi
 12'b101100001101: begin out_real=16'b1110100010110001; out_imag=16'b1100010001100101; end // in_theta = 1.381348 pi
 12'b101100001110: begin out_real=16'b1110100011001001; out_imag=16'b1100010001011100; end // in_theta = 1.381836 pi
 12'b101100001111: begin out_real=16'b1110100011100000; out_imag=16'b1100010001010011; end // in_theta = 1.382324 pi
 12'b101100010000: begin out_real=16'b1110100011110111; out_imag=16'b1100010001001010; end // in_theta = 1.382813 pi
 12'b101100010001: begin out_real=16'b1110100100001111; out_imag=16'b1100010001000001; end // in_theta = 1.383301 pi
 12'b101100010010: begin out_real=16'b1110100100100110; out_imag=16'b1100010000111000; end // in_theta = 1.383789 pi
 12'b101100010011: begin out_real=16'b1110100100111110; out_imag=16'b1100010000101111; end // in_theta = 1.384277 pi
 12'b101100010100: begin out_real=16'b1110100101010101; out_imag=16'b1100010000100110; end // in_theta = 1.384766 pi
 12'b101100010101: begin out_real=16'b1110100101101101; out_imag=16'b1100010000011101; end // in_theta = 1.385254 pi
 12'b101100010110: begin out_real=16'b1110100110000100; out_imag=16'b1100010000010100; end // in_theta = 1.385742 pi
 12'b101100010111: begin out_real=16'b1110100110011100; out_imag=16'b1100010000001011; end // in_theta = 1.386230 pi
 12'b101100011000: begin out_real=16'b1110100110110100; out_imag=16'b1100010000000011; end // in_theta = 1.386719 pi
 12'b101100011001: begin out_real=16'b1110100111001011; out_imag=16'b1100001111111010; end // in_theta = 1.387207 pi
 12'b101100011010: begin out_real=16'b1110100111100011; out_imag=16'b1100001111110001; end // in_theta = 1.387695 pi
 12'b101100011011: begin out_real=16'b1110100111111010; out_imag=16'b1100001111101001; end // in_theta = 1.388184 pi
 12'b101100011100: begin out_real=16'b1110101000010010; out_imag=16'b1100001111100000; end // in_theta = 1.388672 pi
 12'b101100011101: begin out_real=16'b1110101000101001; out_imag=16'b1100001111010111; end // in_theta = 1.389160 pi
 12'b101100011110: begin out_real=16'b1110101001000001; out_imag=16'b1100001111001111; end // in_theta = 1.389648 pi
 12'b101100011111: begin out_real=16'b1110101001011001; out_imag=16'b1100001111000110; end // in_theta = 1.390137 pi
 12'b101100100000: begin out_real=16'b1110101001110000; out_imag=16'b1100001110111110; end // in_theta = 1.390625 pi
 12'b101100100001: begin out_real=16'b1110101010001000; out_imag=16'b1100001110110101; end // in_theta = 1.391113 pi
 12'b101100100010: begin out_real=16'b1110101010100000; out_imag=16'b1100001110101101; end // in_theta = 1.391602 pi
 12'b101100100011: begin out_real=16'b1110101010110111; out_imag=16'b1100001110100101; end // in_theta = 1.392090 pi
 12'b101100100100: begin out_real=16'b1110101011001111; out_imag=16'b1100001110011100; end // in_theta = 1.392578 pi
 12'b101100100101: begin out_real=16'b1110101011100111; out_imag=16'b1100001110010100; end // in_theta = 1.393066 pi
 12'b101100100110: begin out_real=16'b1110101011111111; out_imag=16'b1100001110001100; end // in_theta = 1.393555 pi
 12'b101100100111: begin out_real=16'b1110101100010110; out_imag=16'b1100001110000011; end // in_theta = 1.394043 pi
 12'b101100101000: begin out_real=16'b1110101100101110; out_imag=16'b1100001101111011; end // in_theta = 1.394531 pi
 12'b101100101001: begin out_real=16'b1110101101000110; out_imag=16'b1100001101110011; end // in_theta = 1.395020 pi
 12'b101100101010: begin out_real=16'b1110101101011110; out_imag=16'b1100001101101011; end // in_theta = 1.395508 pi
 12'b101100101011: begin out_real=16'b1110101101110101; out_imag=16'b1100001101100011; end // in_theta = 1.395996 pi
 12'b101100101100: begin out_real=16'b1110101110001101; out_imag=16'b1100001101011011; end // in_theta = 1.396484 pi
 12'b101100101101: begin out_real=16'b1110101110100101; out_imag=16'b1100001101010011; end // in_theta = 1.396973 pi
 12'b101100101110: begin out_real=16'b1110101110111101; out_imag=16'b1100001101001011; end // in_theta = 1.397461 pi
 12'b101100101111: begin out_real=16'b1110101111010101; out_imag=16'b1100001101000011; end // in_theta = 1.397949 pi
 12'b101100110000: begin out_real=16'b1110101111101101; out_imag=16'b1100001100111011; end // in_theta = 1.398438 pi
 12'b101100110001: begin out_real=16'b1110110000000101; out_imag=16'b1100001100110011; end // in_theta = 1.398926 pi
 12'b101100110010: begin out_real=16'b1110110000011100; out_imag=16'b1100001100101011; end // in_theta = 1.399414 pi
 12'b101100110011: begin out_real=16'b1110110000110100; out_imag=16'b1100001100100011; end // in_theta = 1.399902 pi
 12'b101100110100: begin out_real=16'b1110110001001100; out_imag=16'b1100001100011100; end // in_theta = 1.400391 pi
 12'b101100110101: begin out_real=16'b1110110001100100; out_imag=16'b1100001100010100; end // in_theta = 1.400879 pi
 12'b101100110110: begin out_real=16'b1110110001111100; out_imag=16'b1100001100001100; end // in_theta = 1.401367 pi
 12'b101100110111: begin out_real=16'b1110110010010100; out_imag=16'b1100001100000101; end // in_theta = 1.401855 pi
 12'b101100111000: begin out_real=16'b1110110010101100; out_imag=16'b1100001011111101; end // in_theta = 1.402344 pi
 12'b101100111001: begin out_real=16'b1110110011000100; out_imag=16'b1100001011110101; end // in_theta = 1.402832 pi
 12'b101100111010: begin out_real=16'b1110110011011100; out_imag=16'b1100001011101110; end // in_theta = 1.403320 pi
 12'b101100111011: begin out_real=16'b1110110011110100; out_imag=16'b1100001011100110; end // in_theta = 1.403809 pi
 12'b101100111100: begin out_real=16'b1110110100001100; out_imag=16'b1100001011011111; end // in_theta = 1.404297 pi
 12'b101100111101: begin out_real=16'b1110110100100100; out_imag=16'b1100001011011000; end // in_theta = 1.404785 pi
 12'b101100111110: begin out_real=16'b1110110100111100; out_imag=16'b1100001011010000; end // in_theta = 1.405273 pi
 12'b101100111111: begin out_real=16'b1110110101010100; out_imag=16'b1100001011001001; end // in_theta = 1.405762 pi
 12'b101101000000: begin out_real=16'b1110110101101100; out_imag=16'b1100001011000001; end // in_theta = 1.406250 pi
 12'b101101000001: begin out_real=16'b1110110110000100; out_imag=16'b1100001010111010; end // in_theta = 1.406738 pi
 12'b101101000010: begin out_real=16'b1110110110011100; out_imag=16'b1100001010110011; end // in_theta = 1.407227 pi
 12'b101101000011: begin out_real=16'b1110110110110100; out_imag=16'b1100001010101100; end // in_theta = 1.407715 pi
 12'b101101000100: begin out_real=16'b1110110111001100; out_imag=16'b1100001010100101; end // in_theta = 1.408203 pi
 12'b101101000101: begin out_real=16'b1110110111100100; out_imag=16'b1100001010011101; end // in_theta = 1.408691 pi
 12'b101101000110: begin out_real=16'b1110110111111100; out_imag=16'b1100001010010110; end // in_theta = 1.409180 pi
 12'b101101000111: begin out_real=16'b1110111000010101; out_imag=16'b1100001010001111; end // in_theta = 1.409668 pi
 12'b101101001000: begin out_real=16'b1110111000101101; out_imag=16'b1100001010001000; end // in_theta = 1.410156 pi
 12'b101101001001: begin out_real=16'b1110111001000101; out_imag=16'b1100001010000001; end // in_theta = 1.410645 pi
 12'b101101001010: begin out_real=16'b1110111001011101; out_imag=16'b1100001001111010; end // in_theta = 1.411133 pi
 12'b101101001011: begin out_real=16'b1110111001110101; out_imag=16'b1100001001110011; end // in_theta = 1.411621 pi
 12'b101101001100: begin out_real=16'b1110111010001101; out_imag=16'b1100001001101101; end // in_theta = 1.412109 pi
 12'b101101001101: begin out_real=16'b1110111010100110; out_imag=16'b1100001001100110; end // in_theta = 1.412598 pi
 12'b101101001110: begin out_real=16'b1110111010111110; out_imag=16'b1100001001011111; end // in_theta = 1.413086 pi
 12'b101101001111: begin out_real=16'b1110111011010110; out_imag=16'b1100001001011000; end // in_theta = 1.413574 pi
 12'b101101010000: begin out_real=16'b1110111011101110; out_imag=16'b1100001001010001; end // in_theta = 1.414063 pi
 12'b101101010001: begin out_real=16'b1110111100000110; out_imag=16'b1100001001001011; end // in_theta = 1.414551 pi
 12'b101101010010: begin out_real=16'b1110111100011111; out_imag=16'b1100001001000100; end // in_theta = 1.415039 pi
 12'b101101010011: begin out_real=16'b1110111100110111; out_imag=16'b1100001000111110; end // in_theta = 1.415527 pi
 12'b101101010100: begin out_real=16'b1110111101001111; out_imag=16'b1100001000110111; end // in_theta = 1.416016 pi
 12'b101101010101: begin out_real=16'b1110111101100111; out_imag=16'b1100001000110000; end // in_theta = 1.416504 pi
 12'b101101010110: begin out_real=16'b1110111110000000; out_imag=16'b1100001000101010; end // in_theta = 1.416992 pi
 12'b101101010111: begin out_real=16'b1110111110011000; out_imag=16'b1100001000100011; end // in_theta = 1.417480 pi
 12'b101101011000: begin out_real=16'b1110111110110000; out_imag=16'b1100001000011101; end // in_theta = 1.417969 pi
 12'b101101011001: begin out_real=16'b1110111111001001; out_imag=16'b1100001000010111; end // in_theta = 1.418457 pi
 12'b101101011010: begin out_real=16'b1110111111100001; out_imag=16'b1100001000010000; end // in_theta = 1.418945 pi
 12'b101101011011: begin out_real=16'b1110111111111001; out_imag=16'b1100001000001010; end // in_theta = 1.419434 pi
 12'b101101011100: begin out_real=16'b1111000000010010; out_imag=16'b1100001000000100; end // in_theta = 1.419922 pi
 12'b101101011101: begin out_real=16'b1111000000101010; out_imag=16'b1100000111111101; end // in_theta = 1.420410 pi
 12'b101101011110: begin out_real=16'b1111000001000010; out_imag=16'b1100000111110111; end // in_theta = 1.420898 pi
 12'b101101011111: begin out_real=16'b1111000001011011; out_imag=16'b1100000111110001; end // in_theta = 1.421387 pi
 12'b101101100000: begin out_real=16'b1111000001110011; out_imag=16'b1100000111101011; end // in_theta = 1.421875 pi
 12'b101101100001: begin out_real=16'b1111000010001011; out_imag=16'b1100000111100101; end // in_theta = 1.422363 pi
 12'b101101100010: begin out_real=16'b1111000010100100; out_imag=16'b1100000111011111; end // in_theta = 1.422852 pi
 12'b101101100011: begin out_real=16'b1111000010111100; out_imag=16'b1100000111011001; end // in_theta = 1.423340 pi
 12'b101101100100: begin out_real=16'b1111000011010101; out_imag=16'b1100000111010011; end // in_theta = 1.423828 pi
 12'b101101100101: begin out_real=16'b1111000011101101; out_imag=16'b1100000111001101; end // in_theta = 1.424316 pi
 12'b101101100110: begin out_real=16'b1111000100000101; out_imag=16'b1100000111000111; end // in_theta = 1.424805 pi
 12'b101101100111: begin out_real=16'b1111000100011110; out_imag=16'b1100000111000001; end // in_theta = 1.425293 pi
 12'b101101101000: begin out_real=16'b1111000100110110; out_imag=16'b1100000110111011; end // in_theta = 1.425781 pi
 12'b101101101001: begin out_real=16'b1111000101001111; out_imag=16'b1100000110110110; end // in_theta = 1.426270 pi
 12'b101101101010: begin out_real=16'b1111000101100111; out_imag=16'b1100000110110000; end // in_theta = 1.426758 pi
 12'b101101101011: begin out_real=16'b1111000110000000; out_imag=16'b1100000110101010; end // in_theta = 1.427246 pi
 12'b101101101100: begin out_real=16'b1111000110011000; out_imag=16'b1100000110100100; end // in_theta = 1.427734 pi
 12'b101101101101: begin out_real=16'b1111000110110001; out_imag=16'b1100000110011111; end // in_theta = 1.428223 pi
 12'b101101101110: begin out_real=16'b1111000111001001; out_imag=16'b1100000110011001; end // in_theta = 1.428711 pi
 12'b101101101111: begin out_real=16'b1111000111100010; out_imag=16'b1100000110010100; end // in_theta = 1.429199 pi
 12'b101101110000: begin out_real=16'b1111000111111010; out_imag=16'b1100000110001110; end // in_theta = 1.429688 pi
 12'b101101110001: begin out_real=16'b1111001000010011; out_imag=16'b1100000110001001; end // in_theta = 1.430176 pi
 12'b101101110010: begin out_real=16'b1111001000101011; out_imag=16'b1100000110000011; end // in_theta = 1.430664 pi
 12'b101101110011: begin out_real=16'b1111001001000100; out_imag=16'b1100000101111110; end // in_theta = 1.431152 pi
 12'b101101110100: begin out_real=16'b1111001001011100; out_imag=16'b1100000101111000; end // in_theta = 1.431641 pi
 12'b101101110101: begin out_real=16'b1111001001110101; out_imag=16'b1100000101110011; end // in_theta = 1.432129 pi
 12'b101101110110: begin out_real=16'b1111001010001110; out_imag=16'b1100000101101110; end // in_theta = 1.432617 pi
 12'b101101110111: begin out_real=16'b1111001010100110; out_imag=16'b1100000101101000; end // in_theta = 1.433105 pi
 12'b101101111000: begin out_real=16'b1111001010111111; out_imag=16'b1100000101100011; end // in_theta = 1.433594 pi
 12'b101101111001: begin out_real=16'b1111001011010111; out_imag=16'b1100000101011110; end // in_theta = 1.434082 pi
 12'b101101111010: begin out_real=16'b1111001011110000; out_imag=16'b1100000101011001; end // in_theta = 1.434570 pi
 12'b101101111011: begin out_real=16'b1111001100001000; out_imag=16'b1100000101010100; end // in_theta = 1.435059 pi
 12'b101101111100: begin out_real=16'b1111001100100001; out_imag=16'b1100000101001111; end // in_theta = 1.435547 pi
 12'b101101111101: begin out_real=16'b1111001100111010; out_imag=16'b1100000101001010; end // in_theta = 1.436035 pi
 12'b101101111110: begin out_real=16'b1111001101010010; out_imag=16'b1100000101000101; end // in_theta = 1.436523 pi
 12'b101101111111: begin out_real=16'b1111001101101011; out_imag=16'b1100000101000000; end // in_theta = 1.437012 pi
 12'b101110000000: begin out_real=16'b1111001110000100; out_imag=16'b1100000100111011; end // in_theta = 1.437500 pi
 12'b101110000001: begin out_real=16'b1111001110011100; out_imag=16'b1100000100110110; end // in_theta = 1.437988 pi
 12'b101110000010: begin out_real=16'b1111001110110101; out_imag=16'b1100000100110001; end // in_theta = 1.438477 pi
 12'b101110000011: begin out_real=16'b1111001111001110; out_imag=16'b1100000100101100; end // in_theta = 1.438965 pi
 12'b101110000100: begin out_real=16'b1111001111100110; out_imag=16'b1100000100101000; end // in_theta = 1.439453 pi
 12'b101110000101: begin out_real=16'b1111001111111111; out_imag=16'b1100000100100011; end // in_theta = 1.439941 pi
 12'b101110000110: begin out_real=16'b1111010000011000; out_imag=16'b1100000100011110; end // in_theta = 1.440430 pi
 12'b101110000111: begin out_real=16'b1111010000110000; out_imag=16'b1100000100011001; end // in_theta = 1.440918 pi
 12'b101110001000: begin out_real=16'b1111010001001001; out_imag=16'b1100000100010101; end // in_theta = 1.441406 pi
 12'b101110001001: begin out_real=16'b1111010001100010; out_imag=16'b1100000100010000; end // in_theta = 1.441895 pi
 12'b101110001010: begin out_real=16'b1111010001111011; out_imag=16'b1100000100001100; end // in_theta = 1.442383 pi
 12'b101110001011: begin out_real=16'b1111010010010011; out_imag=16'b1100000100000111; end // in_theta = 1.442871 pi
 12'b101110001100: begin out_real=16'b1111010010101100; out_imag=16'b1100000100000011; end // in_theta = 1.443359 pi
 12'b101110001101: begin out_real=16'b1111010011000101; out_imag=16'b1100000011111110; end // in_theta = 1.443848 pi
 12'b101110001110: begin out_real=16'b1111010011011101; out_imag=16'b1100000011111010; end // in_theta = 1.444336 pi
 12'b101110001111: begin out_real=16'b1111010011110110; out_imag=16'b1100000011110110; end // in_theta = 1.444824 pi
 12'b101110010000: begin out_real=16'b1111010100001111; out_imag=16'b1100000011110001; end // in_theta = 1.445313 pi
 12'b101110010001: begin out_real=16'b1111010100101000; out_imag=16'b1100000011101101; end // in_theta = 1.445801 pi
 12'b101110010010: begin out_real=16'b1111010101000000; out_imag=16'b1100000011101001; end // in_theta = 1.446289 pi
 12'b101110010011: begin out_real=16'b1111010101011001; out_imag=16'b1100000011100100; end // in_theta = 1.446777 pi
 12'b101110010100: begin out_real=16'b1111010101110010; out_imag=16'b1100000011100000; end // in_theta = 1.447266 pi
 12'b101110010101: begin out_real=16'b1111010110001011; out_imag=16'b1100000011011100; end // in_theta = 1.447754 pi
 12'b101110010110: begin out_real=16'b1111010110100100; out_imag=16'b1100000011011000; end // in_theta = 1.448242 pi
 12'b101110010111: begin out_real=16'b1111010110111100; out_imag=16'b1100000011010100; end // in_theta = 1.448730 pi
 12'b101110011000: begin out_real=16'b1111010111010101; out_imag=16'b1100000011010000; end // in_theta = 1.449219 pi
 12'b101110011001: begin out_real=16'b1111010111101110; out_imag=16'b1100000011001100; end // in_theta = 1.449707 pi
 12'b101110011010: begin out_real=16'b1111011000000111; out_imag=16'b1100000011001000; end // in_theta = 1.450195 pi
 12'b101110011011: begin out_real=16'b1111011000100000; out_imag=16'b1100000011000100; end // in_theta = 1.450684 pi
 12'b101110011100: begin out_real=16'b1111011000111001; out_imag=16'b1100000011000000; end // in_theta = 1.451172 pi
 12'b101110011101: begin out_real=16'b1111011001010001; out_imag=16'b1100000010111101; end // in_theta = 1.451660 pi
 12'b101110011110: begin out_real=16'b1111011001101010; out_imag=16'b1100000010111001; end // in_theta = 1.452148 pi
 12'b101110011111: begin out_real=16'b1111011010000011; out_imag=16'b1100000010110101; end // in_theta = 1.452637 pi
 12'b101110100000: begin out_real=16'b1111011010011100; out_imag=16'b1100000010110001; end // in_theta = 1.453125 pi
 12'b101110100001: begin out_real=16'b1111011010110101; out_imag=16'b1100000010101110; end // in_theta = 1.453613 pi
 12'b101110100010: begin out_real=16'b1111011011001110; out_imag=16'b1100000010101010; end // in_theta = 1.454102 pi
 12'b101110100011: begin out_real=16'b1111011011100111; out_imag=16'b1100000010100110; end // in_theta = 1.454590 pi
 12'b101110100100: begin out_real=16'b1111011011111111; out_imag=16'b1100000010100011; end // in_theta = 1.455078 pi
 12'b101110100101: begin out_real=16'b1111011100011000; out_imag=16'b1100000010011111; end // in_theta = 1.455566 pi
 12'b101110100110: begin out_real=16'b1111011100110001; out_imag=16'b1100000010011100; end // in_theta = 1.456055 pi
 12'b101110100111: begin out_real=16'b1111011101001010; out_imag=16'b1100000010011000; end // in_theta = 1.456543 pi
 12'b101110101000: begin out_real=16'b1111011101100011; out_imag=16'b1100000010010101; end // in_theta = 1.457031 pi
 12'b101110101001: begin out_real=16'b1111011101111100; out_imag=16'b1100000010010010; end // in_theta = 1.457520 pi
 12'b101110101010: begin out_real=16'b1111011110010101; out_imag=16'b1100000010001110; end // in_theta = 1.458008 pi
 12'b101110101011: begin out_real=16'b1111011110101110; out_imag=16'b1100000010001011; end // in_theta = 1.458496 pi
 12'b101110101100: begin out_real=16'b1111011111000111; out_imag=16'b1100000010001000; end // in_theta = 1.458984 pi
 12'b101110101101: begin out_real=16'b1111011111100000; out_imag=16'b1100000010000101; end // in_theta = 1.459473 pi
 12'b101110101110: begin out_real=16'b1111011111111001; out_imag=16'b1100000010000001; end // in_theta = 1.459961 pi
 12'b101110101111: begin out_real=16'b1111100000010001; out_imag=16'b1100000001111110; end // in_theta = 1.460449 pi
 12'b101110110000: begin out_real=16'b1111100000101010; out_imag=16'b1100000001111011; end // in_theta = 1.460938 pi
 12'b101110110001: begin out_real=16'b1111100001000011; out_imag=16'b1100000001111000; end // in_theta = 1.461426 pi
 12'b101110110010: begin out_real=16'b1111100001011100; out_imag=16'b1100000001110101; end // in_theta = 1.461914 pi
 12'b101110110011: begin out_real=16'b1111100001110101; out_imag=16'b1100000001110010; end // in_theta = 1.462402 pi
 12'b101110110100: begin out_real=16'b1111100010001110; out_imag=16'b1100000001101111; end // in_theta = 1.462891 pi
 12'b101110110101: begin out_real=16'b1111100010100111; out_imag=16'b1100000001101100; end // in_theta = 1.463379 pi
 12'b101110110110: begin out_real=16'b1111100011000000; out_imag=16'b1100000001101001; end // in_theta = 1.463867 pi
 12'b101110110111: begin out_real=16'b1111100011011001; out_imag=16'b1100000001100111; end // in_theta = 1.464355 pi
 12'b101110111000: begin out_real=16'b1111100011110010; out_imag=16'b1100000001100100; end // in_theta = 1.464844 pi
 12'b101110111001: begin out_real=16'b1111100100001011; out_imag=16'b1100000001100001; end // in_theta = 1.465332 pi
 12'b101110111010: begin out_real=16'b1111100100100100; out_imag=16'b1100000001011110; end // in_theta = 1.465820 pi
 12'b101110111011: begin out_real=16'b1111100100111101; out_imag=16'b1100000001011100; end // in_theta = 1.466309 pi
 12'b101110111100: begin out_real=16'b1111100101010110; out_imag=16'b1100000001011001; end // in_theta = 1.466797 pi
 12'b101110111101: begin out_real=16'b1111100101101111; out_imag=16'b1100000001010110; end // in_theta = 1.467285 pi
 12'b101110111110: begin out_real=16'b1111100110001000; out_imag=16'b1100000001010100; end // in_theta = 1.467773 pi
 12'b101110111111: begin out_real=16'b1111100110100001; out_imag=16'b1100000001010001; end // in_theta = 1.468262 pi
 12'b101111000000: begin out_real=16'b1111100110111010; out_imag=16'b1100000001001111; end // in_theta = 1.468750 pi
 12'b101111000001: begin out_real=16'b1111100111010011; out_imag=16'b1100000001001100; end // in_theta = 1.469238 pi
 12'b101111000010: begin out_real=16'b1111100111101100; out_imag=16'b1100000001001010; end // in_theta = 1.469727 pi
 12'b101111000011: begin out_real=16'b1111101000000101; out_imag=16'b1100000001001000; end // in_theta = 1.470215 pi
 12'b101111000100: begin out_real=16'b1111101000011110; out_imag=16'b1100000001000101; end // in_theta = 1.470703 pi
 12'b101111000101: begin out_real=16'b1111101000110111; out_imag=16'b1100000001000011; end // in_theta = 1.471191 pi
 12'b101111000110: begin out_real=16'b1111101001010000; out_imag=16'b1100000001000001; end // in_theta = 1.471680 pi
 12'b101111000111: begin out_real=16'b1111101001101001; out_imag=16'b1100000000111111; end // in_theta = 1.472168 pi
 12'b101111001000: begin out_real=16'b1111101010000010; out_imag=16'b1100000000111100; end // in_theta = 1.472656 pi
 12'b101111001001: begin out_real=16'b1111101010011011; out_imag=16'b1100000000111010; end // in_theta = 1.473145 pi
 12'b101111001010: begin out_real=16'b1111101010110100; out_imag=16'b1100000000111000; end // in_theta = 1.473633 pi
 12'b101111001011: begin out_real=16'b1111101011001101; out_imag=16'b1100000000110110; end // in_theta = 1.474121 pi
 12'b101111001100: begin out_real=16'b1111101011100110; out_imag=16'b1100000000110100; end // in_theta = 1.474609 pi
 12'b101111001101: begin out_real=16'b1111101100000000; out_imag=16'b1100000000110010; end // in_theta = 1.475098 pi
 12'b101111001110: begin out_real=16'b1111101100011001; out_imag=16'b1100000000110000; end // in_theta = 1.475586 pi
 12'b101111001111: begin out_real=16'b1111101100110010; out_imag=16'b1100000000101110; end // in_theta = 1.476074 pi
 12'b101111010000: begin out_real=16'b1111101101001011; out_imag=16'b1100000000101100; end // in_theta = 1.476563 pi
 12'b101111010001: begin out_real=16'b1111101101100100; out_imag=16'b1100000000101011; end // in_theta = 1.477051 pi
 12'b101111010010: begin out_real=16'b1111101101111101; out_imag=16'b1100000000101001; end // in_theta = 1.477539 pi
 12'b101111010011: begin out_real=16'b1111101110010110; out_imag=16'b1100000000100111; end // in_theta = 1.478027 pi
 12'b101111010100: begin out_real=16'b1111101110101111; out_imag=16'b1100000000100101; end // in_theta = 1.478516 pi
 12'b101111010101: begin out_real=16'b1111101111001000; out_imag=16'b1100000000100100; end // in_theta = 1.479004 pi
 12'b101111010110: begin out_real=16'b1111101111100001; out_imag=16'b1100000000100010; end // in_theta = 1.479492 pi
 12'b101111010111: begin out_real=16'b1111101111111010; out_imag=16'b1100000000100000; end // in_theta = 1.479980 pi
 12'b101111011000: begin out_real=16'b1111110000010011; out_imag=16'b1100000000011111; end // in_theta = 1.480469 pi
 12'b101111011001: begin out_real=16'b1111110000101100; out_imag=16'b1100000000011101; end // in_theta = 1.480957 pi
 12'b101111011010: begin out_real=16'b1111110001000101; out_imag=16'b1100000000011100; end // in_theta = 1.481445 pi
 12'b101111011011: begin out_real=16'b1111110001011111; out_imag=16'b1100000000011010; end // in_theta = 1.481934 pi
 12'b101111011100: begin out_real=16'b1111110001111000; out_imag=16'b1100000000011001; end // in_theta = 1.482422 pi
 12'b101111011101: begin out_real=16'b1111110010010001; out_imag=16'b1100000000011000; end // in_theta = 1.482910 pi
 12'b101111011110: begin out_real=16'b1111110010101010; out_imag=16'b1100000000010110; end // in_theta = 1.483398 pi
 12'b101111011111: begin out_real=16'b1111110011000011; out_imag=16'b1100000000010101; end // in_theta = 1.483887 pi
 12'b101111100000: begin out_real=16'b1111110011011100; out_imag=16'b1100000000010100; end // in_theta = 1.484375 pi
 12'b101111100001: begin out_real=16'b1111110011110101; out_imag=16'b1100000000010011; end // in_theta = 1.484863 pi
 12'b101111100010: begin out_real=16'b1111110100001110; out_imag=16'b1100000000010001; end // in_theta = 1.485352 pi
 12'b101111100011: begin out_real=16'b1111110100100111; out_imag=16'b1100000000010000; end // in_theta = 1.485840 pi
 12'b101111100100: begin out_real=16'b1111110101000000; out_imag=16'b1100000000001111; end // in_theta = 1.486328 pi
 12'b101111100101: begin out_real=16'b1111110101011010; out_imag=16'b1100000000001110; end // in_theta = 1.486816 pi
 12'b101111100110: begin out_real=16'b1111110101110011; out_imag=16'b1100000000001101; end // in_theta = 1.487305 pi
 12'b101111100111: begin out_real=16'b1111110110001100; out_imag=16'b1100000000001100; end // in_theta = 1.487793 pi
 12'b101111101000: begin out_real=16'b1111110110100101; out_imag=16'b1100000000001011; end // in_theta = 1.488281 pi
 12'b101111101001: begin out_real=16'b1111110110111110; out_imag=16'b1100000000001010; end // in_theta = 1.488770 pi
 12'b101111101010: begin out_real=16'b1111110111010111; out_imag=16'b1100000000001001; end // in_theta = 1.489258 pi
 12'b101111101011: begin out_real=16'b1111110111110000; out_imag=16'b1100000000001001; end // in_theta = 1.489746 pi
 12'b101111101100: begin out_real=16'b1111111000001001; out_imag=16'b1100000000001000; end // in_theta = 1.490234 pi
 12'b101111101101: begin out_real=16'b1111111000100011; out_imag=16'b1100000000000111; end // in_theta = 1.490723 pi
 12'b101111101110: begin out_real=16'b1111111000111100; out_imag=16'b1100000000000110; end // in_theta = 1.491211 pi
 12'b101111101111: begin out_real=16'b1111111001010101; out_imag=16'b1100000000000110; end // in_theta = 1.491699 pi
 12'b101111110000: begin out_real=16'b1111111001101110; out_imag=16'b1100000000000101; end // in_theta = 1.492188 pi
 12'b101111110001: begin out_real=16'b1111111010000111; out_imag=16'b1100000000000100; end // in_theta = 1.492676 pi
 12'b101111110010: begin out_real=16'b1111111010100000; out_imag=16'b1100000000000100; end // in_theta = 1.493164 pi
 12'b101111110011: begin out_real=16'b1111111010111001; out_imag=16'b1100000000000011; end // in_theta = 1.493652 pi
 12'b101111110100: begin out_real=16'b1111111011010010; out_imag=16'b1100000000000011; end // in_theta = 1.494141 pi
 12'b101111110101: begin out_real=16'b1111111011101100; out_imag=16'b1100000000000010; end // in_theta = 1.494629 pi
 12'b101111110110: begin out_real=16'b1111111100000101; out_imag=16'b1100000000000010; end // in_theta = 1.495117 pi
 12'b101111110111: begin out_real=16'b1111111100011110; out_imag=16'b1100000000000010; end // in_theta = 1.495605 pi
 12'b101111111000: begin out_real=16'b1111111100110111; out_imag=16'b1100000000000001; end // in_theta = 1.496094 pi
 12'b101111111001: begin out_real=16'b1111111101010000; out_imag=16'b1100000000000001; end // in_theta = 1.496582 pi
 12'b101111111010: begin out_real=16'b1111111101101001; out_imag=16'b1100000000000001; end // in_theta = 1.497070 pi
 12'b101111111011: begin out_real=16'b1111111110000010; out_imag=16'b1100000000000000; end // in_theta = 1.497559 pi
 12'b101111111100: begin out_real=16'b1111111110011011; out_imag=16'b1100000000000000; end // in_theta = 1.498047 pi
 12'b101111111101: begin out_real=16'b1111111110110101; out_imag=16'b1100000000000000; end // in_theta = 1.498535 pi
 12'b101111111110: begin out_real=16'b1111111111001110; out_imag=16'b1100000000000000; end // in_theta = 1.499023 pi
 12'b101111111111: begin out_real=16'b1111111111100111; out_imag=16'b1100000000000000; end // in_theta = 1.499512 pi
 12'b110000000000: begin out_real=16'b0000000000000000; out_imag=16'b1100000000000000; end // in_theta = 1.500000 pi
 12'b110000000001: begin out_real=16'b0000000000011001; out_imag=16'b1100000000000000; end // in_theta = 1.500488 pi
 12'b110000000010: begin out_real=16'b0000000000110010; out_imag=16'b1100000000000000; end // in_theta = 1.500977 pi
 12'b110000000011: begin out_real=16'b0000000001001011; out_imag=16'b1100000000000000; end // in_theta = 1.501465 pi
 12'b110000000100: begin out_real=16'b0000000001100101; out_imag=16'b1100000000000000; end // in_theta = 1.501953 pi
 12'b110000000101: begin out_real=16'b0000000001111110; out_imag=16'b1100000000000000; end // in_theta = 1.502441 pi
 12'b110000000110: begin out_real=16'b0000000010010111; out_imag=16'b1100000000000001; end // in_theta = 1.502930 pi
 12'b110000000111: begin out_real=16'b0000000010110000; out_imag=16'b1100000000000001; end // in_theta = 1.503418 pi
 12'b110000001000: begin out_real=16'b0000000011001001; out_imag=16'b1100000000000001; end // in_theta = 1.503906 pi
 12'b110000001001: begin out_real=16'b0000000011100010; out_imag=16'b1100000000000010; end // in_theta = 1.504395 pi
 12'b110000001010: begin out_real=16'b0000000011111011; out_imag=16'b1100000000000010; end // in_theta = 1.504883 pi
 12'b110000001011: begin out_real=16'b0000000100010100; out_imag=16'b1100000000000010; end // in_theta = 1.505371 pi
 12'b110000001100: begin out_real=16'b0000000100101110; out_imag=16'b1100000000000011; end // in_theta = 1.505859 pi
 12'b110000001101: begin out_real=16'b0000000101000111; out_imag=16'b1100000000000011; end // in_theta = 1.506348 pi
 12'b110000001110: begin out_real=16'b0000000101100000; out_imag=16'b1100000000000100; end // in_theta = 1.506836 pi
 12'b110000001111: begin out_real=16'b0000000101111001; out_imag=16'b1100000000000100; end // in_theta = 1.507324 pi
 12'b110000010000: begin out_real=16'b0000000110010010; out_imag=16'b1100000000000101; end // in_theta = 1.507813 pi
 12'b110000010001: begin out_real=16'b0000000110101011; out_imag=16'b1100000000000110; end // in_theta = 1.508301 pi
 12'b110000010010: begin out_real=16'b0000000111000100; out_imag=16'b1100000000000110; end // in_theta = 1.508789 pi
 12'b110000010011: begin out_real=16'b0000000111011101; out_imag=16'b1100000000000111; end // in_theta = 1.509277 pi
 12'b110000010100: begin out_real=16'b0000000111110111; out_imag=16'b1100000000001000; end // in_theta = 1.509766 pi
 12'b110000010101: begin out_real=16'b0000001000010000; out_imag=16'b1100000000001001; end // in_theta = 1.510254 pi
 12'b110000010110: begin out_real=16'b0000001000101001; out_imag=16'b1100000000001001; end // in_theta = 1.510742 pi
 12'b110000010111: begin out_real=16'b0000001001000010; out_imag=16'b1100000000001010; end // in_theta = 1.511230 pi
 12'b110000011000: begin out_real=16'b0000001001011011; out_imag=16'b1100000000001011; end // in_theta = 1.511719 pi
 12'b110000011001: begin out_real=16'b0000001001110100; out_imag=16'b1100000000001100; end // in_theta = 1.512207 pi
 12'b110000011010: begin out_real=16'b0000001010001101; out_imag=16'b1100000000001101; end // in_theta = 1.512695 pi
 12'b110000011011: begin out_real=16'b0000001010100110; out_imag=16'b1100000000001110; end // in_theta = 1.513184 pi
 12'b110000011100: begin out_real=16'b0000001011000000; out_imag=16'b1100000000001111; end // in_theta = 1.513672 pi
 12'b110000011101: begin out_real=16'b0000001011011001; out_imag=16'b1100000000010000; end // in_theta = 1.514160 pi
 12'b110000011110: begin out_real=16'b0000001011110010; out_imag=16'b1100000000010001; end // in_theta = 1.514648 pi
 12'b110000011111: begin out_real=16'b0000001100001011; out_imag=16'b1100000000010011; end // in_theta = 1.515137 pi
 12'b110000100000: begin out_real=16'b0000001100100100; out_imag=16'b1100000000010100; end // in_theta = 1.515625 pi
 12'b110000100001: begin out_real=16'b0000001100111101; out_imag=16'b1100000000010101; end // in_theta = 1.516113 pi
 12'b110000100010: begin out_real=16'b0000001101010110; out_imag=16'b1100000000010110; end // in_theta = 1.516602 pi
 12'b110000100011: begin out_real=16'b0000001101101111; out_imag=16'b1100000000011000; end // in_theta = 1.517090 pi
 12'b110000100100: begin out_real=16'b0000001110001000; out_imag=16'b1100000000011001; end // in_theta = 1.517578 pi
 12'b110000100101: begin out_real=16'b0000001110100001; out_imag=16'b1100000000011010; end // in_theta = 1.518066 pi
 12'b110000100110: begin out_real=16'b0000001110111011; out_imag=16'b1100000000011100; end // in_theta = 1.518555 pi
 12'b110000100111: begin out_real=16'b0000001111010100; out_imag=16'b1100000000011101; end // in_theta = 1.519043 pi
 12'b110000101000: begin out_real=16'b0000001111101101; out_imag=16'b1100000000011111; end // in_theta = 1.519531 pi
 12'b110000101001: begin out_real=16'b0000010000000110; out_imag=16'b1100000000100000; end // in_theta = 1.520020 pi
 12'b110000101010: begin out_real=16'b0000010000011111; out_imag=16'b1100000000100010; end // in_theta = 1.520508 pi
 12'b110000101011: begin out_real=16'b0000010000111000; out_imag=16'b1100000000100100; end // in_theta = 1.520996 pi
 12'b110000101100: begin out_real=16'b0000010001010001; out_imag=16'b1100000000100101; end // in_theta = 1.521484 pi
 12'b110000101101: begin out_real=16'b0000010001101010; out_imag=16'b1100000000100111; end // in_theta = 1.521973 pi
 12'b110000101110: begin out_real=16'b0000010010000011; out_imag=16'b1100000000101001; end // in_theta = 1.522461 pi
 12'b110000101111: begin out_real=16'b0000010010011100; out_imag=16'b1100000000101011; end // in_theta = 1.522949 pi
 12'b110000110000: begin out_real=16'b0000010010110101; out_imag=16'b1100000000101100; end // in_theta = 1.523438 pi
 12'b110000110001: begin out_real=16'b0000010011001110; out_imag=16'b1100000000101110; end // in_theta = 1.523926 pi
 12'b110000110010: begin out_real=16'b0000010011100111; out_imag=16'b1100000000110000; end // in_theta = 1.524414 pi
 12'b110000110011: begin out_real=16'b0000010100000000; out_imag=16'b1100000000110010; end // in_theta = 1.524902 pi
 12'b110000110100: begin out_real=16'b0000010100011010; out_imag=16'b1100000000110100; end // in_theta = 1.525391 pi
 12'b110000110101: begin out_real=16'b0000010100110011; out_imag=16'b1100000000110110; end // in_theta = 1.525879 pi
 12'b110000110110: begin out_real=16'b0000010101001100; out_imag=16'b1100000000111000; end // in_theta = 1.526367 pi
 12'b110000110111: begin out_real=16'b0000010101100101; out_imag=16'b1100000000111010; end // in_theta = 1.526855 pi
 12'b110000111000: begin out_real=16'b0000010101111110; out_imag=16'b1100000000111100; end // in_theta = 1.527344 pi
 12'b110000111001: begin out_real=16'b0000010110010111; out_imag=16'b1100000000111111; end // in_theta = 1.527832 pi
 12'b110000111010: begin out_real=16'b0000010110110000; out_imag=16'b1100000001000001; end // in_theta = 1.528320 pi
 12'b110000111011: begin out_real=16'b0000010111001001; out_imag=16'b1100000001000011; end // in_theta = 1.528809 pi
 12'b110000111100: begin out_real=16'b0000010111100010; out_imag=16'b1100000001000101; end // in_theta = 1.529297 pi
 12'b110000111101: begin out_real=16'b0000010111111011; out_imag=16'b1100000001001000; end // in_theta = 1.529785 pi
 12'b110000111110: begin out_real=16'b0000011000010100; out_imag=16'b1100000001001010; end // in_theta = 1.530273 pi
 12'b110000111111: begin out_real=16'b0000011000101101; out_imag=16'b1100000001001100; end // in_theta = 1.530762 pi
 12'b110001000000: begin out_real=16'b0000011001000110; out_imag=16'b1100000001001111; end // in_theta = 1.531250 pi
 12'b110001000001: begin out_real=16'b0000011001011111; out_imag=16'b1100000001010001; end // in_theta = 1.531738 pi
 12'b110001000010: begin out_real=16'b0000011001111000; out_imag=16'b1100000001010100; end // in_theta = 1.532227 pi
 12'b110001000011: begin out_real=16'b0000011010010001; out_imag=16'b1100000001010110; end // in_theta = 1.532715 pi
 12'b110001000100: begin out_real=16'b0000011010101010; out_imag=16'b1100000001011001; end // in_theta = 1.533203 pi
 12'b110001000101: begin out_real=16'b0000011011000011; out_imag=16'b1100000001011100; end // in_theta = 1.533691 pi
 12'b110001000110: begin out_real=16'b0000011011011100; out_imag=16'b1100000001011110; end // in_theta = 1.534180 pi
 12'b110001000111: begin out_real=16'b0000011011110101; out_imag=16'b1100000001100001; end // in_theta = 1.534668 pi
 12'b110001001000: begin out_real=16'b0000011100001110; out_imag=16'b1100000001100100; end // in_theta = 1.535156 pi
 12'b110001001001: begin out_real=16'b0000011100100111; out_imag=16'b1100000001100111; end // in_theta = 1.535645 pi
 12'b110001001010: begin out_real=16'b0000011101000000; out_imag=16'b1100000001101001; end // in_theta = 1.536133 pi
 12'b110001001011: begin out_real=16'b0000011101011001; out_imag=16'b1100000001101100; end // in_theta = 1.536621 pi
 12'b110001001100: begin out_real=16'b0000011101110010; out_imag=16'b1100000001101111; end // in_theta = 1.537109 pi
 12'b110001001101: begin out_real=16'b0000011110001011; out_imag=16'b1100000001110010; end // in_theta = 1.537598 pi
 12'b110001001110: begin out_real=16'b0000011110100100; out_imag=16'b1100000001110101; end // in_theta = 1.538086 pi
 12'b110001001111: begin out_real=16'b0000011110111101; out_imag=16'b1100000001111000; end // in_theta = 1.538574 pi
 12'b110001010000: begin out_real=16'b0000011111010110; out_imag=16'b1100000001111011; end // in_theta = 1.539062 pi
 12'b110001010001: begin out_real=16'b0000011111101111; out_imag=16'b1100000001111110; end // in_theta = 1.539551 pi
 12'b110001010010: begin out_real=16'b0000100000000111; out_imag=16'b1100000010000001; end // in_theta = 1.540039 pi
 12'b110001010011: begin out_real=16'b0000100000100000; out_imag=16'b1100000010000101; end // in_theta = 1.540527 pi
 12'b110001010100: begin out_real=16'b0000100000111001; out_imag=16'b1100000010001000; end // in_theta = 1.541016 pi
 12'b110001010101: begin out_real=16'b0000100001010010; out_imag=16'b1100000010001011; end // in_theta = 1.541504 pi
 12'b110001010110: begin out_real=16'b0000100001101011; out_imag=16'b1100000010001110; end // in_theta = 1.541992 pi
 12'b110001010111: begin out_real=16'b0000100010000100; out_imag=16'b1100000010010010; end // in_theta = 1.542480 pi
 12'b110001011000: begin out_real=16'b0000100010011101; out_imag=16'b1100000010010101; end // in_theta = 1.542969 pi
 12'b110001011001: begin out_real=16'b0000100010110110; out_imag=16'b1100000010011000; end // in_theta = 1.543457 pi
 12'b110001011010: begin out_real=16'b0000100011001111; out_imag=16'b1100000010011100; end // in_theta = 1.543945 pi
 12'b110001011011: begin out_real=16'b0000100011101000; out_imag=16'b1100000010011111; end // in_theta = 1.544434 pi
 12'b110001011100: begin out_real=16'b0000100100000001; out_imag=16'b1100000010100011; end // in_theta = 1.544922 pi
 12'b110001011101: begin out_real=16'b0000100100011001; out_imag=16'b1100000010100110; end // in_theta = 1.545410 pi
 12'b110001011110: begin out_real=16'b0000100100110010; out_imag=16'b1100000010101010; end // in_theta = 1.545898 pi
 12'b110001011111: begin out_real=16'b0000100101001011; out_imag=16'b1100000010101110; end // in_theta = 1.546387 pi
 12'b110001100000: begin out_real=16'b0000100101100100; out_imag=16'b1100000010110001; end // in_theta = 1.546875 pi
 12'b110001100001: begin out_real=16'b0000100101111101; out_imag=16'b1100000010110101; end // in_theta = 1.547363 pi
 12'b110001100010: begin out_real=16'b0000100110010110; out_imag=16'b1100000010111001; end // in_theta = 1.547852 pi
 12'b110001100011: begin out_real=16'b0000100110101111; out_imag=16'b1100000010111101; end // in_theta = 1.548340 pi
 12'b110001100100: begin out_real=16'b0000100111000111; out_imag=16'b1100000011000000; end // in_theta = 1.548828 pi
 12'b110001100101: begin out_real=16'b0000100111100000; out_imag=16'b1100000011000100; end // in_theta = 1.549316 pi
 12'b110001100110: begin out_real=16'b0000100111111001; out_imag=16'b1100000011001000; end // in_theta = 1.549805 pi
 12'b110001100111: begin out_real=16'b0000101000010010; out_imag=16'b1100000011001100; end // in_theta = 1.550293 pi
 12'b110001101000: begin out_real=16'b0000101000101011; out_imag=16'b1100000011010000; end // in_theta = 1.550781 pi
 12'b110001101001: begin out_real=16'b0000101001000100; out_imag=16'b1100000011010100; end // in_theta = 1.551270 pi
 12'b110001101010: begin out_real=16'b0000101001011100; out_imag=16'b1100000011011000; end // in_theta = 1.551758 pi
 12'b110001101011: begin out_real=16'b0000101001110101; out_imag=16'b1100000011011100; end // in_theta = 1.552246 pi
 12'b110001101100: begin out_real=16'b0000101010001110; out_imag=16'b1100000011100000; end // in_theta = 1.552734 pi
 12'b110001101101: begin out_real=16'b0000101010100111; out_imag=16'b1100000011100100; end // in_theta = 1.553223 pi
 12'b110001101110: begin out_real=16'b0000101011000000; out_imag=16'b1100000011101001; end // in_theta = 1.553711 pi
 12'b110001101111: begin out_real=16'b0000101011011000; out_imag=16'b1100000011101101; end // in_theta = 1.554199 pi
 12'b110001110000: begin out_real=16'b0000101011110001; out_imag=16'b1100000011110001; end // in_theta = 1.554688 pi
 12'b110001110001: begin out_real=16'b0000101100001010; out_imag=16'b1100000011110110; end // in_theta = 1.555176 pi
 12'b110001110010: begin out_real=16'b0000101100100011; out_imag=16'b1100000011111010; end // in_theta = 1.555664 pi
 12'b110001110011: begin out_real=16'b0000101100111011; out_imag=16'b1100000011111110; end // in_theta = 1.556152 pi
 12'b110001110100: begin out_real=16'b0000101101010100; out_imag=16'b1100000100000011; end // in_theta = 1.556641 pi
 12'b110001110101: begin out_real=16'b0000101101101101; out_imag=16'b1100000100000111; end // in_theta = 1.557129 pi
 12'b110001110110: begin out_real=16'b0000101110000101; out_imag=16'b1100000100001100; end // in_theta = 1.557617 pi
 12'b110001110111: begin out_real=16'b0000101110011110; out_imag=16'b1100000100010000; end // in_theta = 1.558105 pi
 12'b110001111000: begin out_real=16'b0000101110110111; out_imag=16'b1100000100010101; end // in_theta = 1.558594 pi
 12'b110001111001: begin out_real=16'b0000101111010000; out_imag=16'b1100000100011001; end // in_theta = 1.559082 pi
 12'b110001111010: begin out_real=16'b0000101111101000; out_imag=16'b1100000100011110; end // in_theta = 1.559570 pi
 12'b110001111011: begin out_real=16'b0000110000000001; out_imag=16'b1100000100100011; end // in_theta = 1.560059 pi
 12'b110001111100: begin out_real=16'b0000110000011010; out_imag=16'b1100000100101000; end // in_theta = 1.560547 pi
 12'b110001111101: begin out_real=16'b0000110000110010; out_imag=16'b1100000100101100; end // in_theta = 1.561035 pi
 12'b110001111110: begin out_real=16'b0000110001001011; out_imag=16'b1100000100110001; end // in_theta = 1.561523 pi
 12'b110001111111: begin out_real=16'b0000110001100100; out_imag=16'b1100000100110110; end // in_theta = 1.562012 pi
 12'b110010000000: begin out_real=16'b0000110001111100; out_imag=16'b1100000100111011; end // in_theta = 1.562500 pi
 12'b110010000001: begin out_real=16'b0000110010010101; out_imag=16'b1100000101000000; end // in_theta = 1.562988 pi
 12'b110010000010: begin out_real=16'b0000110010101110; out_imag=16'b1100000101000101; end // in_theta = 1.563477 pi
 12'b110010000011: begin out_real=16'b0000110011000110; out_imag=16'b1100000101001010; end // in_theta = 1.563965 pi
 12'b110010000100: begin out_real=16'b0000110011011111; out_imag=16'b1100000101001111; end // in_theta = 1.564453 pi
 12'b110010000101: begin out_real=16'b0000110011111000; out_imag=16'b1100000101010100; end // in_theta = 1.564941 pi
 12'b110010000110: begin out_real=16'b0000110100010000; out_imag=16'b1100000101011001; end // in_theta = 1.565430 pi
 12'b110010000111: begin out_real=16'b0000110100101001; out_imag=16'b1100000101011110; end // in_theta = 1.565918 pi
 12'b110010001000: begin out_real=16'b0000110101000001; out_imag=16'b1100000101100011; end // in_theta = 1.566406 pi
 12'b110010001001: begin out_real=16'b0000110101011010; out_imag=16'b1100000101101000; end // in_theta = 1.566895 pi
 12'b110010001010: begin out_real=16'b0000110101110010; out_imag=16'b1100000101101110; end // in_theta = 1.567383 pi
 12'b110010001011: begin out_real=16'b0000110110001011; out_imag=16'b1100000101110011; end // in_theta = 1.567871 pi
 12'b110010001100: begin out_real=16'b0000110110100100; out_imag=16'b1100000101111000; end // in_theta = 1.568359 pi
 12'b110010001101: begin out_real=16'b0000110110111100; out_imag=16'b1100000101111110; end // in_theta = 1.568848 pi
 12'b110010001110: begin out_real=16'b0000110111010101; out_imag=16'b1100000110000011; end // in_theta = 1.569336 pi
 12'b110010001111: begin out_real=16'b0000110111101101; out_imag=16'b1100000110001001; end // in_theta = 1.569824 pi
 12'b110010010000: begin out_real=16'b0000111000000110; out_imag=16'b1100000110001110; end // in_theta = 1.570313 pi
 12'b110010010001: begin out_real=16'b0000111000011110; out_imag=16'b1100000110010100; end // in_theta = 1.570801 pi
 12'b110010010010: begin out_real=16'b0000111000110111; out_imag=16'b1100000110011001; end // in_theta = 1.571289 pi
 12'b110010010011: begin out_real=16'b0000111001001111; out_imag=16'b1100000110011111; end // in_theta = 1.571777 pi
 12'b110010010100: begin out_real=16'b0000111001101000; out_imag=16'b1100000110100100; end // in_theta = 1.572266 pi
 12'b110010010101: begin out_real=16'b0000111010000000; out_imag=16'b1100000110101010; end // in_theta = 1.572754 pi
 12'b110010010110: begin out_real=16'b0000111010011001; out_imag=16'b1100000110110000; end // in_theta = 1.573242 pi
 12'b110010010111: begin out_real=16'b0000111010110001; out_imag=16'b1100000110110110; end // in_theta = 1.573730 pi
 12'b110010011000: begin out_real=16'b0000111011001010; out_imag=16'b1100000110111011; end // in_theta = 1.574219 pi
 12'b110010011001: begin out_real=16'b0000111011100010; out_imag=16'b1100000111000001; end // in_theta = 1.574707 pi
 12'b110010011010: begin out_real=16'b0000111011111011; out_imag=16'b1100000111000111; end // in_theta = 1.575195 pi
 12'b110010011011: begin out_real=16'b0000111100010011; out_imag=16'b1100000111001101; end // in_theta = 1.575684 pi
 12'b110010011100: begin out_real=16'b0000111100101011; out_imag=16'b1100000111010011; end // in_theta = 1.576172 pi
 12'b110010011101: begin out_real=16'b0000111101000100; out_imag=16'b1100000111011001; end // in_theta = 1.576660 pi
 12'b110010011110: begin out_real=16'b0000111101011100; out_imag=16'b1100000111011111; end // in_theta = 1.577148 pi
 12'b110010011111: begin out_real=16'b0000111101110101; out_imag=16'b1100000111100101; end // in_theta = 1.577637 pi
 12'b110010100000: begin out_real=16'b0000111110001101; out_imag=16'b1100000111101011; end // in_theta = 1.578125 pi
 12'b110010100001: begin out_real=16'b0000111110100101; out_imag=16'b1100000111110001; end // in_theta = 1.578613 pi
 12'b110010100010: begin out_real=16'b0000111110111110; out_imag=16'b1100000111110111; end // in_theta = 1.579102 pi
 12'b110010100011: begin out_real=16'b0000111111010110; out_imag=16'b1100000111111101; end // in_theta = 1.579590 pi
 12'b110010100100: begin out_real=16'b0000111111101110; out_imag=16'b1100001000000100; end // in_theta = 1.580078 pi
 12'b110010100101: begin out_real=16'b0001000000000111; out_imag=16'b1100001000001010; end // in_theta = 1.580566 pi
 12'b110010100110: begin out_real=16'b0001000000011111; out_imag=16'b1100001000010000; end // in_theta = 1.581055 pi
 12'b110010100111: begin out_real=16'b0001000000110111; out_imag=16'b1100001000010111; end // in_theta = 1.581543 pi
 12'b110010101000: begin out_real=16'b0001000001010000; out_imag=16'b1100001000011101; end // in_theta = 1.582031 pi
 12'b110010101001: begin out_real=16'b0001000001101000; out_imag=16'b1100001000100011; end // in_theta = 1.582520 pi
 12'b110010101010: begin out_real=16'b0001000010000000; out_imag=16'b1100001000101010; end // in_theta = 1.583008 pi
 12'b110010101011: begin out_real=16'b0001000010011001; out_imag=16'b1100001000110000; end // in_theta = 1.583496 pi
 12'b110010101100: begin out_real=16'b0001000010110001; out_imag=16'b1100001000110111; end // in_theta = 1.583984 pi
 12'b110010101101: begin out_real=16'b0001000011001001; out_imag=16'b1100001000111110; end // in_theta = 1.584473 pi
 12'b110010101110: begin out_real=16'b0001000011100001; out_imag=16'b1100001001000100; end // in_theta = 1.584961 pi
 12'b110010101111: begin out_real=16'b0001000011111010; out_imag=16'b1100001001001011; end // in_theta = 1.585449 pi
 12'b110010110000: begin out_real=16'b0001000100010010; out_imag=16'b1100001001010001; end // in_theta = 1.585938 pi
 12'b110010110001: begin out_real=16'b0001000100101010; out_imag=16'b1100001001011000; end // in_theta = 1.586426 pi
 12'b110010110010: begin out_real=16'b0001000101000010; out_imag=16'b1100001001011111; end // in_theta = 1.586914 pi
 12'b110010110011: begin out_real=16'b0001000101011010; out_imag=16'b1100001001100110; end // in_theta = 1.587402 pi
 12'b110010110100: begin out_real=16'b0001000101110011; out_imag=16'b1100001001101101; end // in_theta = 1.587891 pi
 12'b110010110101: begin out_real=16'b0001000110001011; out_imag=16'b1100001001110011; end // in_theta = 1.588379 pi
 12'b110010110110: begin out_real=16'b0001000110100011; out_imag=16'b1100001001111010; end // in_theta = 1.588867 pi
 12'b110010110111: begin out_real=16'b0001000110111011; out_imag=16'b1100001010000001; end // in_theta = 1.589355 pi
 12'b110010111000: begin out_real=16'b0001000111010011; out_imag=16'b1100001010001000; end // in_theta = 1.589844 pi
 12'b110010111001: begin out_real=16'b0001000111101011; out_imag=16'b1100001010001111; end // in_theta = 1.590332 pi
 12'b110010111010: begin out_real=16'b0001001000000100; out_imag=16'b1100001010010110; end // in_theta = 1.590820 pi
 12'b110010111011: begin out_real=16'b0001001000011100; out_imag=16'b1100001010011101; end // in_theta = 1.591309 pi
 12'b110010111100: begin out_real=16'b0001001000110100; out_imag=16'b1100001010100101; end // in_theta = 1.591797 pi
 12'b110010111101: begin out_real=16'b0001001001001100; out_imag=16'b1100001010101100; end // in_theta = 1.592285 pi
 12'b110010111110: begin out_real=16'b0001001001100100; out_imag=16'b1100001010110011; end // in_theta = 1.592773 pi
 12'b110010111111: begin out_real=16'b0001001001111100; out_imag=16'b1100001010111010; end // in_theta = 1.593262 pi
 12'b110011000000: begin out_real=16'b0001001010010100; out_imag=16'b1100001011000001; end // in_theta = 1.593750 pi
 12'b110011000001: begin out_real=16'b0001001010101100; out_imag=16'b1100001011001001; end // in_theta = 1.594238 pi
 12'b110011000010: begin out_real=16'b0001001011000100; out_imag=16'b1100001011010000; end // in_theta = 1.594727 pi
 12'b110011000011: begin out_real=16'b0001001011011100; out_imag=16'b1100001011011000; end // in_theta = 1.595215 pi
 12'b110011000100: begin out_real=16'b0001001011110100; out_imag=16'b1100001011011111; end // in_theta = 1.595703 pi
 12'b110011000101: begin out_real=16'b0001001100001100; out_imag=16'b1100001011100110; end // in_theta = 1.596191 pi
 12'b110011000110: begin out_real=16'b0001001100100100; out_imag=16'b1100001011101110; end // in_theta = 1.596680 pi
 12'b110011000111: begin out_real=16'b0001001100111100; out_imag=16'b1100001011110101; end // in_theta = 1.597168 pi
 12'b110011001000: begin out_real=16'b0001001101010100; out_imag=16'b1100001011111101; end // in_theta = 1.597656 pi
 12'b110011001001: begin out_real=16'b0001001101101100; out_imag=16'b1100001100000101; end // in_theta = 1.598145 pi
 12'b110011001010: begin out_real=16'b0001001110000100; out_imag=16'b1100001100001100; end // in_theta = 1.598633 pi
 12'b110011001011: begin out_real=16'b0001001110011100; out_imag=16'b1100001100010100; end // in_theta = 1.599121 pi
 12'b110011001100: begin out_real=16'b0001001110110100; out_imag=16'b1100001100011100; end // in_theta = 1.599609 pi
 12'b110011001101: begin out_real=16'b0001001111001100; out_imag=16'b1100001100100011; end // in_theta = 1.600098 pi
 12'b110011001110: begin out_real=16'b0001001111100100; out_imag=16'b1100001100101011; end // in_theta = 1.600586 pi
 12'b110011001111: begin out_real=16'b0001001111111011; out_imag=16'b1100001100110011; end // in_theta = 1.601074 pi
 12'b110011010000: begin out_real=16'b0001010000010011; out_imag=16'b1100001100111011; end // in_theta = 1.601563 pi
 12'b110011010001: begin out_real=16'b0001010000101011; out_imag=16'b1100001101000011; end // in_theta = 1.602051 pi
 12'b110011010010: begin out_real=16'b0001010001000011; out_imag=16'b1100001101001011; end // in_theta = 1.602539 pi
 12'b110011010011: begin out_real=16'b0001010001011011; out_imag=16'b1100001101010011; end // in_theta = 1.603027 pi
 12'b110011010100: begin out_real=16'b0001010001110011; out_imag=16'b1100001101011011; end // in_theta = 1.603516 pi
 12'b110011010101: begin out_real=16'b0001010010001011; out_imag=16'b1100001101100011; end // in_theta = 1.604004 pi
 12'b110011010110: begin out_real=16'b0001010010100010; out_imag=16'b1100001101101011; end // in_theta = 1.604492 pi
 12'b110011010111: begin out_real=16'b0001010010111010; out_imag=16'b1100001101110011; end // in_theta = 1.604980 pi
 12'b110011011000: begin out_real=16'b0001010011010010; out_imag=16'b1100001101111011; end // in_theta = 1.605469 pi
 12'b110011011001: begin out_real=16'b0001010011101010; out_imag=16'b1100001110000011; end // in_theta = 1.605957 pi
 12'b110011011010: begin out_real=16'b0001010100000001; out_imag=16'b1100001110001100; end // in_theta = 1.606445 pi
 12'b110011011011: begin out_real=16'b0001010100011001; out_imag=16'b1100001110010100; end // in_theta = 1.606934 pi
 12'b110011011100: begin out_real=16'b0001010100110001; out_imag=16'b1100001110011100; end // in_theta = 1.607422 pi
 12'b110011011101: begin out_real=16'b0001010101001001; out_imag=16'b1100001110100101; end // in_theta = 1.607910 pi
 12'b110011011110: begin out_real=16'b0001010101100000; out_imag=16'b1100001110101101; end // in_theta = 1.608398 pi
 12'b110011011111: begin out_real=16'b0001010101111000; out_imag=16'b1100001110110101; end // in_theta = 1.608887 pi
 12'b110011100000: begin out_real=16'b0001010110010000; out_imag=16'b1100001110111110; end // in_theta = 1.609375 pi
 12'b110011100001: begin out_real=16'b0001010110100111; out_imag=16'b1100001111000110; end // in_theta = 1.609863 pi
 12'b110011100010: begin out_real=16'b0001010110111111; out_imag=16'b1100001111001111; end // in_theta = 1.610352 pi
 12'b110011100011: begin out_real=16'b0001010111010111; out_imag=16'b1100001111010111; end // in_theta = 1.610840 pi
 12'b110011100100: begin out_real=16'b0001010111101110; out_imag=16'b1100001111100000; end // in_theta = 1.611328 pi
 12'b110011100101: begin out_real=16'b0001011000000110; out_imag=16'b1100001111101001; end // in_theta = 1.611816 pi
 12'b110011100110: begin out_real=16'b0001011000011101; out_imag=16'b1100001111110001; end // in_theta = 1.612305 pi
 12'b110011100111: begin out_real=16'b0001011000110101; out_imag=16'b1100001111111010; end // in_theta = 1.612793 pi
 12'b110011101000: begin out_real=16'b0001011001001100; out_imag=16'b1100010000000011; end // in_theta = 1.613281 pi
 12'b110011101001: begin out_real=16'b0001011001100100; out_imag=16'b1100010000001011; end // in_theta = 1.613770 pi
 12'b110011101010: begin out_real=16'b0001011001111100; out_imag=16'b1100010000010100; end // in_theta = 1.614258 pi
 12'b110011101011: begin out_real=16'b0001011010010011; out_imag=16'b1100010000011101; end // in_theta = 1.614746 pi
 12'b110011101100: begin out_real=16'b0001011010101011; out_imag=16'b1100010000100110; end // in_theta = 1.615234 pi
 12'b110011101101: begin out_real=16'b0001011011000010; out_imag=16'b1100010000101111; end // in_theta = 1.615723 pi
 12'b110011101110: begin out_real=16'b0001011011011010; out_imag=16'b1100010000111000; end // in_theta = 1.616211 pi
 12'b110011101111: begin out_real=16'b0001011011110001; out_imag=16'b1100010001000001; end // in_theta = 1.616699 pi
 12'b110011110000: begin out_real=16'b0001011100001001; out_imag=16'b1100010001001010; end // in_theta = 1.617187 pi
 12'b110011110001: begin out_real=16'b0001011100100000; out_imag=16'b1100010001010011; end // in_theta = 1.617676 pi
 12'b110011110010: begin out_real=16'b0001011100110111; out_imag=16'b1100010001011100; end // in_theta = 1.618164 pi
 12'b110011110011: begin out_real=16'b0001011101001111; out_imag=16'b1100010001100101; end // in_theta = 1.618652 pi
 12'b110011110100: begin out_real=16'b0001011101100110; out_imag=16'b1100010001101110; end // in_theta = 1.619141 pi
 12'b110011110101: begin out_real=16'b0001011101111110; out_imag=16'b1100010001111000; end // in_theta = 1.619629 pi
 12'b110011110110: begin out_real=16'b0001011110010101; out_imag=16'b1100010010000001; end // in_theta = 1.620117 pi
 12'b110011110111: begin out_real=16'b0001011110101100; out_imag=16'b1100010010001010; end // in_theta = 1.620605 pi
 12'b110011111000: begin out_real=16'b0001011111000100; out_imag=16'b1100010010010011; end // in_theta = 1.621094 pi
 12'b110011111001: begin out_real=16'b0001011111011011; out_imag=16'b1100010010011101; end // in_theta = 1.621582 pi
 12'b110011111010: begin out_real=16'b0001011111110010; out_imag=16'b1100010010100110; end // in_theta = 1.622070 pi
 12'b110011111011: begin out_real=16'b0001100000001010; out_imag=16'b1100010010110000; end // in_theta = 1.622559 pi
 12'b110011111100: begin out_real=16'b0001100000100001; out_imag=16'b1100010010111001; end // in_theta = 1.623047 pi
 12'b110011111101: begin out_real=16'b0001100000111000; out_imag=16'b1100010011000010; end // in_theta = 1.623535 pi
 12'b110011111110: begin out_real=16'b0001100001001111; out_imag=16'b1100010011001100; end // in_theta = 1.624023 pi
 12'b110011111111: begin out_real=16'b0001100001100111; out_imag=16'b1100010011010110; end // in_theta = 1.624512 pi
 12'b110100000000: begin out_real=16'b0001100001111110; out_imag=16'b1100010011011111; end // in_theta = 1.625000 pi
 12'b110100000001: begin out_real=16'b0001100010010101; out_imag=16'b1100010011101001; end // in_theta = 1.625488 pi
 12'b110100000010: begin out_real=16'b0001100010101100; out_imag=16'b1100010011110010; end // in_theta = 1.625977 pi
 12'b110100000011: begin out_real=16'b0001100011000011; out_imag=16'b1100010011111100; end // in_theta = 1.626465 pi
 12'b110100000100: begin out_real=16'b0001100011011011; out_imag=16'b1100010100000110; end // in_theta = 1.626953 pi
 12'b110100000101: begin out_real=16'b0001100011110010; out_imag=16'b1100010100010000; end // in_theta = 1.627441 pi
 12'b110100000110: begin out_real=16'b0001100100001001; out_imag=16'b1100010100011010; end // in_theta = 1.627930 pi
 12'b110100000111: begin out_real=16'b0001100100100000; out_imag=16'b1100010100100011; end // in_theta = 1.628418 pi
 12'b110100001000: begin out_real=16'b0001100100110111; out_imag=16'b1100010100101101; end // in_theta = 1.628906 pi
 12'b110100001001: begin out_real=16'b0001100101001110; out_imag=16'b1100010100110111; end // in_theta = 1.629395 pi
 12'b110100001010: begin out_real=16'b0001100101100101; out_imag=16'b1100010101000001; end // in_theta = 1.629883 pi
 12'b110100001011: begin out_real=16'b0001100101111100; out_imag=16'b1100010101001011; end // in_theta = 1.630371 pi
 12'b110100001100: begin out_real=16'b0001100110010011; out_imag=16'b1100010101010101; end // in_theta = 1.630859 pi
 12'b110100001101: begin out_real=16'b0001100110101010; out_imag=16'b1100010101011111; end // in_theta = 1.631348 pi
 12'b110100001110: begin out_real=16'b0001100111000001; out_imag=16'b1100010101101001; end // in_theta = 1.631836 pi
 12'b110100001111: begin out_real=16'b0001100111011000; out_imag=16'b1100010101110011; end // in_theta = 1.632324 pi
 12'b110100010000: begin out_real=16'b0001100111101111; out_imag=16'b1100010101111110; end // in_theta = 1.632813 pi
 12'b110100010001: begin out_real=16'b0001101000000110; out_imag=16'b1100010110001000; end // in_theta = 1.633301 pi
 12'b110100010010: begin out_real=16'b0001101000011101; out_imag=16'b1100010110010010; end // in_theta = 1.633789 pi
 12'b110100010011: begin out_real=16'b0001101000110100; out_imag=16'b1100010110011100; end // in_theta = 1.634277 pi
 12'b110100010100: begin out_real=16'b0001101001001011; out_imag=16'b1100010110100111; end // in_theta = 1.634766 pi
 12'b110100010101: begin out_real=16'b0001101001100010; out_imag=16'b1100010110110001; end // in_theta = 1.635254 pi
 12'b110100010110: begin out_real=16'b0001101001111001; out_imag=16'b1100010110111011; end // in_theta = 1.635742 pi
 12'b110100010111: begin out_real=16'b0001101010010000; out_imag=16'b1100010111000110; end // in_theta = 1.636230 pi
 12'b110100011000: begin out_real=16'b0001101010100111; out_imag=16'b1100010111010000; end // in_theta = 1.636719 pi
 12'b110100011001: begin out_real=16'b0001101010111110; out_imag=16'b1100010111011011; end // in_theta = 1.637207 pi
 12'b110100011010: begin out_real=16'b0001101011010100; out_imag=16'b1100010111100101; end // in_theta = 1.637695 pi
 12'b110100011011: begin out_real=16'b0001101011101011; out_imag=16'b1100010111110000; end // in_theta = 1.638184 pi
 12'b110100011100: begin out_real=16'b0001101100000010; out_imag=16'b1100010111111010; end // in_theta = 1.638672 pi
 12'b110100011101: begin out_real=16'b0001101100011001; out_imag=16'b1100011000000101; end // in_theta = 1.639160 pi
 12'b110100011110: begin out_real=16'b0001101100110000; out_imag=16'b1100011000010000; end // in_theta = 1.639648 pi
 12'b110100011111: begin out_real=16'b0001101101000110; out_imag=16'b1100011000011010; end // in_theta = 1.640137 pi
 12'b110100100000: begin out_real=16'b0001101101011101; out_imag=16'b1100011000100101; end // in_theta = 1.640625 pi
 12'b110100100001: begin out_real=16'b0001101101110100; out_imag=16'b1100011000110000; end // in_theta = 1.641113 pi
 12'b110100100010: begin out_real=16'b0001101110001010; out_imag=16'b1100011000111011; end // in_theta = 1.641602 pi
 12'b110100100011: begin out_real=16'b0001101110100001; out_imag=16'b1100011001000101; end // in_theta = 1.642090 pi
 12'b110100100100: begin out_real=16'b0001101110111000; out_imag=16'b1100011001010000; end // in_theta = 1.642578 pi
 12'b110100100101: begin out_real=16'b0001101111001110; out_imag=16'b1100011001011011; end // in_theta = 1.643066 pi
 12'b110100100110: begin out_real=16'b0001101111100101; out_imag=16'b1100011001100110; end // in_theta = 1.643555 pi
 12'b110100100111: begin out_real=16'b0001101111111100; out_imag=16'b1100011001110001; end // in_theta = 1.644043 pi
 12'b110100101000: begin out_real=16'b0001110000010010; out_imag=16'b1100011001111100; end // in_theta = 1.644531 pi
 12'b110100101001: begin out_real=16'b0001110000101001; out_imag=16'b1100011010000111; end // in_theta = 1.645020 pi
 12'b110100101010: begin out_real=16'b0001110000111111; out_imag=16'b1100011010010010; end // in_theta = 1.645508 pi
 12'b110100101011: begin out_real=16'b0001110001010110; out_imag=16'b1100011010011101; end // in_theta = 1.645996 pi
 12'b110100101100: begin out_real=16'b0001110001101100; out_imag=16'b1100011010101000; end // in_theta = 1.646484 pi
 12'b110100101101: begin out_real=16'b0001110010000011; out_imag=16'b1100011010110100; end // in_theta = 1.646973 pi
 12'b110100101110: begin out_real=16'b0001110010011001; out_imag=16'b1100011010111111; end // in_theta = 1.647461 pi
 12'b110100101111: begin out_real=16'b0001110010110000; out_imag=16'b1100011011001010; end // in_theta = 1.647949 pi
 12'b110100110000: begin out_real=16'b0001110011000110; out_imag=16'b1100011011010101; end // in_theta = 1.648438 pi
 12'b110100110001: begin out_real=16'b0001110011011101; out_imag=16'b1100011011100001; end // in_theta = 1.648926 pi
 12'b110100110010: begin out_real=16'b0001110011110011; out_imag=16'b1100011011101100; end // in_theta = 1.649414 pi
 12'b110100110011: begin out_real=16'b0001110100001010; out_imag=16'b1100011011110111; end // in_theta = 1.649902 pi
 12'b110100110100: begin out_real=16'b0001110100100000; out_imag=16'b1100011100000011; end // in_theta = 1.650391 pi
 12'b110100110101: begin out_real=16'b0001110100110110; out_imag=16'b1100011100001110; end // in_theta = 1.650879 pi
 12'b110100110110: begin out_real=16'b0001110101001101; out_imag=16'b1100011100011010; end // in_theta = 1.651367 pi
 12'b110100110111: begin out_real=16'b0001110101100011; out_imag=16'b1100011100100101; end // in_theta = 1.651855 pi
 12'b110100111000: begin out_real=16'b0001110101111001; out_imag=16'b1100011100110001; end // in_theta = 1.652344 pi
 12'b110100111001: begin out_real=16'b0001110110010000; out_imag=16'b1100011100111101; end // in_theta = 1.652832 pi
 12'b110100111010: begin out_real=16'b0001110110100110; out_imag=16'b1100011101001000; end // in_theta = 1.653320 pi
 12'b110100111011: begin out_real=16'b0001110110111100; out_imag=16'b1100011101010100; end // in_theta = 1.653809 pi
 12'b110100111100: begin out_real=16'b0001110111010011; out_imag=16'b1100011101011111; end // in_theta = 1.654297 pi
 12'b110100111101: begin out_real=16'b0001110111101001; out_imag=16'b1100011101101011; end // in_theta = 1.654785 pi
 12'b110100111110: begin out_real=16'b0001110111111111; out_imag=16'b1100011101110111; end // in_theta = 1.655273 pi
 12'b110100111111: begin out_real=16'b0001111000010101; out_imag=16'b1100011110000011; end // in_theta = 1.655762 pi
 12'b110101000000: begin out_real=16'b0001111000101011; out_imag=16'b1100011110001111; end // in_theta = 1.656250 pi
 12'b110101000001: begin out_real=16'b0001111001000010; out_imag=16'b1100011110011010; end // in_theta = 1.656738 pi
 12'b110101000010: begin out_real=16'b0001111001011000; out_imag=16'b1100011110100110; end // in_theta = 1.657227 pi
 12'b110101000011: begin out_real=16'b0001111001101110; out_imag=16'b1100011110110010; end // in_theta = 1.657715 pi
 12'b110101000100: begin out_real=16'b0001111010000100; out_imag=16'b1100011110111110; end // in_theta = 1.658203 pi
 12'b110101000101: begin out_real=16'b0001111010011010; out_imag=16'b1100011111001010; end // in_theta = 1.658691 pi
 12'b110101000110: begin out_real=16'b0001111010110000; out_imag=16'b1100011111010110; end // in_theta = 1.659180 pi
 12'b110101000111: begin out_real=16'b0001111011000110; out_imag=16'b1100011111100010; end // in_theta = 1.659668 pi
 12'b110101001000: begin out_real=16'b0001111011011100; out_imag=16'b1100011111101110; end // in_theta = 1.660156 pi
 12'b110101001001: begin out_real=16'b0001111011110010; out_imag=16'b1100011111111011; end // in_theta = 1.660645 pi
 12'b110101001010: begin out_real=16'b0001111100001000; out_imag=16'b1100100000000111; end // in_theta = 1.661133 pi
 12'b110101001011: begin out_real=16'b0001111100011110; out_imag=16'b1100100000010011; end // in_theta = 1.661621 pi
 12'b110101001100: begin out_real=16'b0001111100110100; out_imag=16'b1100100000011111; end // in_theta = 1.662109 pi
 12'b110101001101: begin out_real=16'b0001111101001010; out_imag=16'b1100100000101011; end // in_theta = 1.662598 pi
 12'b110101001110: begin out_real=16'b0001111101100000; out_imag=16'b1100100000111000; end // in_theta = 1.663086 pi
 12'b110101001111: begin out_real=16'b0001111101110110; out_imag=16'b1100100001000100; end // in_theta = 1.663574 pi
 12'b110101010000: begin out_real=16'b0001111110001100; out_imag=16'b1100100001010000; end // in_theta = 1.664063 pi
 12'b110101010001: begin out_real=16'b0001111110100010; out_imag=16'b1100100001011101; end // in_theta = 1.664551 pi
 12'b110101010010: begin out_real=16'b0001111110110111; out_imag=16'b1100100001101001; end // in_theta = 1.665039 pi
 12'b110101010011: begin out_real=16'b0001111111001101; out_imag=16'b1100100001110110; end // in_theta = 1.665527 pi
 12'b110101010100: begin out_real=16'b0001111111100011; out_imag=16'b1100100010000010; end // in_theta = 1.666016 pi
 12'b110101010101: begin out_real=16'b0001111111111001; out_imag=16'b1100100010001111; end // in_theta = 1.666504 pi
 12'b110101010110: begin out_real=16'b0010000000001111; out_imag=16'b1100100010011011; end // in_theta = 1.666992 pi
 12'b110101010111: begin out_real=16'b0010000000100100; out_imag=16'b1100100010101000; end // in_theta = 1.667480 pi
 12'b110101011000: begin out_real=16'b0010000000111010; out_imag=16'b1100100010110101; end // in_theta = 1.667969 pi
 12'b110101011001: begin out_real=16'b0010000001010000; out_imag=16'b1100100011000001; end // in_theta = 1.668457 pi
 12'b110101011010: begin out_real=16'b0010000001100101; out_imag=16'b1100100011001110; end // in_theta = 1.668945 pi
 12'b110101011011: begin out_real=16'b0010000001111011; out_imag=16'b1100100011011011; end // in_theta = 1.669434 pi
 12'b110101011100: begin out_real=16'b0010000010010001; out_imag=16'b1100100011101000; end // in_theta = 1.669922 pi
 12'b110101011101: begin out_real=16'b0010000010100110; out_imag=16'b1100100011110100; end // in_theta = 1.670410 pi
 12'b110101011110: begin out_real=16'b0010000010111100; out_imag=16'b1100100100000001; end // in_theta = 1.670898 pi
 12'b110101011111: begin out_real=16'b0010000011010001; out_imag=16'b1100100100001110; end // in_theta = 1.671387 pi
 12'b110101100000: begin out_real=16'b0010000011100111; out_imag=16'b1100100100011011; end // in_theta = 1.671875 pi
 12'b110101100001: begin out_real=16'b0010000011111101; out_imag=16'b1100100100101000; end // in_theta = 1.672363 pi
 12'b110101100010: begin out_real=16'b0010000100010010; out_imag=16'b1100100100110101; end // in_theta = 1.672852 pi
 12'b110101100011: begin out_real=16'b0010000100101000; out_imag=16'b1100100101000010; end // in_theta = 1.673340 pi
 12'b110101100100: begin out_real=16'b0010000100111101; out_imag=16'b1100100101001111; end // in_theta = 1.673828 pi
 12'b110101100101: begin out_real=16'b0010000101010011; out_imag=16'b1100100101011100; end // in_theta = 1.674316 pi
 12'b110101100110: begin out_real=16'b0010000101101000; out_imag=16'b1100100101101001; end // in_theta = 1.674805 pi
 12'b110101100111: begin out_real=16'b0010000101111101; out_imag=16'b1100100101110110; end // in_theta = 1.675293 pi
 12'b110101101000: begin out_real=16'b0010000110010011; out_imag=16'b1100100110000011; end // in_theta = 1.675781 pi
 12'b110101101001: begin out_real=16'b0010000110101000; out_imag=16'b1100100110010001; end // in_theta = 1.676270 pi
 12'b110101101010: begin out_real=16'b0010000110111110; out_imag=16'b1100100110011110; end // in_theta = 1.676758 pi
 12'b110101101011: begin out_real=16'b0010000111010011; out_imag=16'b1100100110101011; end // in_theta = 1.677246 pi
 12'b110101101100: begin out_real=16'b0010000111101000; out_imag=16'b1100100110111000; end // in_theta = 1.677734 pi
 12'b110101101101: begin out_real=16'b0010000111111110; out_imag=16'b1100100111000110; end // in_theta = 1.678223 pi
 12'b110101101110: begin out_real=16'b0010001000010011; out_imag=16'b1100100111010011; end // in_theta = 1.678711 pi
 12'b110101101111: begin out_real=16'b0010001000101000; out_imag=16'b1100100111100000; end // in_theta = 1.679199 pi
 12'b110101110000: begin out_real=16'b0010001000111101; out_imag=16'b1100100111101110; end // in_theta = 1.679688 pi
 12'b110101110001: begin out_real=16'b0010001001010011; out_imag=16'b1100100111111011; end // in_theta = 1.680176 pi
 12'b110101110010: begin out_real=16'b0010001001101000; out_imag=16'b1100101000001001; end // in_theta = 1.680664 pi
 12'b110101110011: begin out_real=16'b0010001001111101; out_imag=16'b1100101000010110; end // in_theta = 1.681152 pi
 12'b110101110100: begin out_real=16'b0010001010010010; out_imag=16'b1100101000100100; end // in_theta = 1.681641 pi
 12'b110101110101: begin out_real=16'b0010001010100111; out_imag=16'b1100101000110010; end // in_theta = 1.682129 pi
 12'b110101110110: begin out_real=16'b0010001010111100; out_imag=16'b1100101000111111; end // in_theta = 1.682617 pi
 12'b110101110111: begin out_real=16'b0010001011010010; out_imag=16'b1100101001001101; end // in_theta = 1.683105 pi
 12'b110101111000: begin out_real=16'b0010001011100111; out_imag=16'b1100101001011011; end // in_theta = 1.683594 pi
 12'b110101111001: begin out_real=16'b0010001011111100; out_imag=16'b1100101001101000; end // in_theta = 1.684082 pi
 12'b110101111010: begin out_real=16'b0010001100010001; out_imag=16'b1100101001110110; end // in_theta = 1.684570 pi
 12'b110101111011: begin out_real=16'b0010001100100110; out_imag=16'b1100101010000100; end // in_theta = 1.685059 pi
 12'b110101111100: begin out_real=16'b0010001100111011; out_imag=16'b1100101010010010; end // in_theta = 1.685547 pi
 12'b110101111101: begin out_real=16'b0010001101010000; out_imag=16'b1100101010011111; end // in_theta = 1.686035 pi
 12'b110101111110: begin out_real=16'b0010001101100101; out_imag=16'b1100101010101101; end // in_theta = 1.686523 pi
 12'b110101111111: begin out_real=16'b0010001101111010; out_imag=16'b1100101010111011; end // in_theta = 1.687012 pi
 12'b110110000000: begin out_real=16'b0010001110001110; out_imag=16'b1100101011001001; end // in_theta = 1.687500 pi
 12'b110110000001: begin out_real=16'b0010001110100011; out_imag=16'b1100101011010111; end // in_theta = 1.687988 pi
 12'b110110000010: begin out_real=16'b0010001110111000; out_imag=16'b1100101011100101; end // in_theta = 1.688477 pi
 12'b110110000011: begin out_real=16'b0010001111001101; out_imag=16'b1100101011110011; end // in_theta = 1.688965 pi
 12'b110110000100: begin out_real=16'b0010001111100010; out_imag=16'b1100101100000001; end // in_theta = 1.689453 pi
 12'b110110000101: begin out_real=16'b0010001111110111; out_imag=16'b1100101100001111; end // in_theta = 1.689941 pi
 12'b110110000110: begin out_real=16'b0010010000001011; out_imag=16'b1100101100011110; end // in_theta = 1.690430 pi
 12'b110110000111: begin out_real=16'b0010010000100000; out_imag=16'b1100101100101100; end // in_theta = 1.690918 pi
 12'b110110001000: begin out_real=16'b0010010000110101; out_imag=16'b1100101100111010; end // in_theta = 1.691406 pi
 12'b110110001001: begin out_real=16'b0010010001001010; out_imag=16'b1100101101001000; end // in_theta = 1.691895 pi
 12'b110110001010: begin out_real=16'b0010010001011110; out_imag=16'b1100101101010110; end // in_theta = 1.692383 pi
 12'b110110001011: begin out_real=16'b0010010001110011; out_imag=16'b1100101101100101; end // in_theta = 1.692871 pi
 12'b110110001100: begin out_real=16'b0010010010001000; out_imag=16'b1100101101110011; end // in_theta = 1.693359 pi
 12'b110110001101: begin out_real=16'b0010010010011100; out_imag=16'b1100101110000001; end // in_theta = 1.693848 pi
 12'b110110001110: begin out_real=16'b0010010010110001; out_imag=16'b1100101110010000; end // in_theta = 1.694336 pi
 12'b110110001111: begin out_real=16'b0010010011000101; out_imag=16'b1100101110011110; end // in_theta = 1.694824 pi
 12'b110110010000: begin out_real=16'b0010010011011010; out_imag=16'b1100101110101101; end // in_theta = 1.695313 pi
 12'b110110010001: begin out_real=16'b0010010011101111; out_imag=16'b1100101110111011; end // in_theta = 1.695801 pi
 12'b110110010010: begin out_real=16'b0010010100000011; out_imag=16'b1100101111001010; end // in_theta = 1.696289 pi
 12'b110110010011: begin out_real=16'b0010010100011000; out_imag=16'b1100101111011000; end // in_theta = 1.696777 pi
 12'b110110010100: begin out_real=16'b0010010100101100; out_imag=16'b1100101111100111; end // in_theta = 1.697266 pi
 12'b110110010101: begin out_real=16'b0010010101000001; out_imag=16'b1100101111110101; end // in_theta = 1.697754 pi
 12'b110110010110: begin out_real=16'b0010010101010101; out_imag=16'b1100110000000100; end // in_theta = 1.698242 pi
 12'b110110010111: begin out_real=16'b0010010101101001; out_imag=16'b1100110000010011; end // in_theta = 1.698730 pi
 12'b110110011000: begin out_real=16'b0010010101111110; out_imag=16'b1100110000100001; end // in_theta = 1.699219 pi
 12'b110110011001: begin out_real=16'b0010010110010010; out_imag=16'b1100110000110000; end // in_theta = 1.699707 pi
 12'b110110011010: begin out_real=16'b0010010110100110; out_imag=16'b1100110000111111; end // in_theta = 1.700195 pi
 12'b110110011011: begin out_real=16'b0010010110111011; out_imag=16'b1100110001001110; end // in_theta = 1.700684 pi
 12'b110110011100: begin out_real=16'b0010010111001111; out_imag=16'b1100110001011101; end // in_theta = 1.701172 pi
 12'b110110011101: begin out_real=16'b0010010111100011; out_imag=16'b1100110001101011; end // in_theta = 1.701660 pi
 12'b110110011110: begin out_real=16'b0010010111111000; out_imag=16'b1100110001111010; end // in_theta = 1.702148 pi
 12'b110110011111: begin out_real=16'b0010011000001100; out_imag=16'b1100110010001001; end // in_theta = 1.702637 pi
 12'b110110100000: begin out_real=16'b0010011000100000; out_imag=16'b1100110010011000; end // in_theta = 1.703125 pi
 12'b110110100001: begin out_real=16'b0010011000110100; out_imag=16'b1100110010100111; end // in_theta = 1.703613 pi
 12'b110110100010: begin out_real=16'b0010011001001000; out_imag=16'b1100110010110110; end // in_theta = 1.704102 pi
 12'b110110100011: begin out_real=16'b0010011001011100; out_imag=16'b1100110011000101; end // in_theta = 1.704590 pi
 12'b110110100100: begin out_real=16'b0010011001110001; out_imag=16'b1100110011010100; end // in_theta = 1.705078 pi
 12'b110110100101: begin out_real=16'b0010011010000101; out_imag=16'b1100110011100011; end // in_theta = 1.705566 pi
 12'b110110100110: begin out_real=16'b0010011010011001; out_imag=16'b1100110011110011; end // in_theta = 1.706055 pi
 12'b110110100111: begin out_real=16'b0010011010101101; out_imag=16'b1100110100000010; end // in_theta = 1.706543 pi
 12'b110110101000: begin out_real=16'b0010011011000001; out_imag=16'b1100110100010001; end // in_theta = 1.707031 pi
 12'b110110101001: begin out_real=16'b0010011011010101; out_imag=16'b1100110100100000; end // in_theta = 1.707520 pi
 12'b110110101010: begin out_real=16'b0010011011101001; out_imag=16'b1100110100110000; end // in_theta = 1.708008 pi
 12'b110110101011: begin out_real=16'b0010011011111101; out_imag=16'b1100110100111111; end // in_theta = 1.708496 pi
 12'b110110101100: begin out_real=16'b0010011100010001; out_imag=16'b1100110101001110; end // in_theta = 1.708984 pi
 12'b110110101101: begin out_real=16'b0010011100100100; out_imag=16'b1100110101011101; end // in_theta = 1.709473 pi
 12'b110110101110: begin out_real=16'b0010011100111000; out_imag=16'b1100110101101101; end // in_theta = 1.709961 pi
 12'b110110101111: begin out_real=16'b0010011101001100; out_imag=16'b1100110101111100; end // in_theta = 1.710449 pi
 12'b110110110000: begin out_real=16'b0010011101100000; out_imag=16'b1100110110001100; end // in_theta = 1.710938 pi
 12'b110110110001: begin out_real=16'b0010011101110100; out_imag=16'b1100110110011011; end // in_theta = 1.711426 pi
 12'b110110110010: begin out_real=16'b0010011110001000; out_imag=16'b1100110110101011; end // in_theta = 1.711914 pi
 12'b110110110011: begin out_real=16'b0010011110011011; out_imag=16'b1100110110111010; end // in_theta = 1.712402 pi
 12'b110110110100: begin out_real=16'b0010011110101111; out_imag=16'b1100110111001010; end // in_theta = 1.712891 pi
 12'b110110110101: begin out_real=16'b0010011111000011; out_imag=16'b1100110111011001; end // in_theta = 1.713379 pi
 12'b110110110110: begin out_real=16'b0010011111010110; out_imag=16'b1100110111101001; end // in_theta = 1.713867 pi
 12'b110110110111: begin out_real=16'b0010011111101010; out_imag=16'b1100110111111001; end // in_theta = 1.714355 pi
 12'b110110111000: begin out_real=16'b0010011111111110; out_imag=16'b1100111000001000; end // in_theta = 1.714844 pi
 12'b110110111001: begin out_real=16'b0010100000010001; out_imag=16'b1100111000011000; end // in_theta = 1.715332 pi
 12'b110110111010: begin out_real=16'b0010100000100101; out_imag=16'b1100111000101000; end // in_theta = 1.715820 pi
 12'b110110111011: begin out_real=16'b0010100000111000; out_imag=16'b1100111000111000; end // in_theta = 1.716309 pi
 12'b110110111100: begin out_real=16'b0010100001001100; out_imag=16'b1100111001000111; end // in_theta = 1.716797 pi
 12'b110110111101: begin out_real=16'b0010100001100000; out_imag=16'b1100111001010111; end // in_theta = 1.717285 pi
 12'b110110111110: begin out_real=16'b0010100001110011; out_imag=16'b1100111001100111; end // in_theta = 1.717773 pi
 12'b110110111111: begin out_real=16'b0010100010000110; out_imag=16'b1100111001110111; end // in_theta = 1.718262 pi
 12'b110111000000: begin out_real=16'b0010100010011010; out_imag=16'b1100111010000111; end // in_theta = 1.718750 pi
 12'b110111000001: begin out_real=16'b0010100010101101; out_imag=16'b1100111010010111; end // in_theta = 1.719238 pi
 12'b110111000010: begin out_real=16'b0010100011000001; out_imag=16'b1100111010100111; end // in_theta = 1.719727 pi
 12'b110111000011: begin out_real=16'b0010100011010100; out_imag=16'b1100111010110111; end // in_theta = 1.720215 pi
 12'b110111000100: begin out_real=16'b0010100011100111; out_imag=16'b1100111011000111; end // in_theta = 1.720703 pi
 12'b110111000101: begin out_real=16'b0010100011111011; out_imag=16'b1100111011010111; end // in_theta = 1.721191 pi
 12'b110111000110: begin out_real=16'b0010100100001110; out_imag=16'b1100111011100111; end // in_theta = 1.721680 pi
 12'b110111000111: begin out_real=16'b0010100100100001; out_imag=16'b1100111011110111; end // in_theta = 1.722168 pi
 12'b110111001000: begin out_real=16'b0010100100110101; out_imag=16'b1100111100000111; end // in_theta = 1.722656 pi
 12'b110111001001: begin out_real=16'b0010100101001000; out_imag=16'b1100111100011000; end // in_theta = 1.723145 pi
 12'b110111001010: begin out_real=16'b0010100101011011; out_imag=16'b1100111100101000; end // in_theta = 1.723633 pi
 12'b110111001011: begin out_real=16'b0010100101101110; out_imag=16'b1100111100111000; end // in_theta = 1.724121 pi
 12'b110111001100: begin out_real=16'b0010100110000001; out_imag=16'b1100111101001000; end // in_theta = 1.724609 pi
 12'b110111001101: begin out_real=16'b0010100110010100; out_imag=16'b1100111101011001; end // in_theta = 1.725098 pi
 12'b110111001110: begin out_real=16'b0010100110100111; out_imag=16'b1100111101101001; end // in_theta = 1.725586 pi
 12'b110111001111: begin out_real=16'b0010100110111011; out_imag=16'b1100111101111001; end // in_theta = 1.726074 pi
 12'b110111010000: begin out_real=16'b0010100111001110; out_imag=16'b1100111110001010; end // in_theta = 1.726563 pi
 12'b110111010001: begin out_real=16'b0010100111100001; out_imag=16'b1100111110011010; end // in_theta = 1.727051 pi
 12'b110111010010: begin out_real=16'b0010100111110100; out_imag=16'b1100111110101011; end // in_theta = 1.727539 pi
 12'b110111010011: begin out_real=16'b0010101000000111; out_imag=16'b1100111110111011; end // in_theta = 1.728027 pi
 12'b110111010100: begin out_real=16'b0010101000011010; out_imag=16'b1100111111001100; end // in_theta = 1.728516 pi
 12'b110111010101: begin out_real=16'b0010101000101100; out_imag=16'b1100111111011100; end // in_theta = 1.729004 pi
 12'b110111010110: begin out_real=16'b0010101000111111; out_imag=16'b1100111111101101; end // in_theta = 1.729492 pi
 12'b110111010111: begin out_real=16'b0010101001010010; out_imag=16'b1100111111111110; end // in_theta = 1.729980 pi
 12'b110111011000: begin out_real=16'b0010101001100101; out_imag=16'b1101000000001110; end // in_theta = 1.730469 pi
 12'b110111011001: begin out_real=16'b0010101001111000; out_imag=16'b1101000000011111; end // in_theta = 1.730957 pi
 12'b110111011010: begin out_real=16'b0010101010001011; out_imag=16'b1101000000110000; end // in_theta = 1.731445 pi
 12'b110111011011: begin out_real=16'b0010101010011101; out_imag=16'b1101000001000000; end // in_theta = 1.731934 pi
 12'b110111011100: begin out_real=16'b0010101010110000; out_imag=16'b1101000001010001; end // in_theta = 1.732422 pi
 12'b110111011101: begin out_real=16'b0010101011000011; out_imag=16'b1101000001100010; end // in_theta = 1.732910 pi
 12'b110111011110: begin out_real=16'b0010101011010110; out_imag=16'b1101000001110011; end // in_theta = 1.733398 pi
 12'b110111011111: begin out_real=16'b0010101011101000; out_imag=16'b1101000010000011; end // in_theta = 1.733887 pi
 12'b110111100000: begin out_real=16'b0010101011111011; out_imag=16'b1101000010010100; end // in_theta = 1.734375 pi
 12'b110111100001: begin out_real=16'b0010101100001101; out_imag=16'b1101000010100101; end // in_theta = 1.734863 pi
 12'b110111100010: begin out_real=16'b0010101100100000; out_imag=16'b1101000010110110; end // in_theta = 1.735352 pi
 12'b110111100011: begin out_real=16'b0010101100110011; out_imag=16'b1101000011000111; end // in_theta = 1.735840 pi
 12'b110111100100: begin out_real=16'b0010101101000101; out_imag=16'b1101000011011000; end // in_theta = 1.736328 pi
 12'b110111100101: begin out_real=16'b0010101101011000; out_imag=16'b1101000011101001; end // in_theta = 1.736816 pi
 12'b110111100110: begin out_real=16'b0010101101101010; out_imag=16'b1101000011111010; end // in_theta = 1.737305 pi
 12'b110111100111: begin out_real=16'b0010101101111101; out_imag=16'b1101000100001011; end // in_theta = 1.737793 pi
 12'b110111101000: begin out_real=16'b0010101110001111; out_imag=16'b1101000100011100; end // in_theta = 1.738281 pi
 12'b110111101001: begin out_real=16'b0010101110100001; out_imag=16'b1101000100101101; end // in_theta = 1.738770 pi
 12'b110111101010: begin out_real=16'b0010101110110100; out_imag=16'b1101000100111110; end // in_theta = 1.739258 pi
 12'b110111101011: begin out_real=16'b0010101111000110; out_imag=16'b1101000101010000; end // in_theta = 1.739746 pi
 12'b110111101100: begin out_real=16'b0010101111011000; out_imag=16'b1101000101100001; end // in_theta = 1.740234 pi
 12'b110111101101: begin out_real=16'b0010101111101011; out_imag=16'b1101000101110010; end // in_theta = 1.740723 pi
 12'b110111101110: begin out_real=16'b0010101111111101; out_imag=16'b1101000110000011; end // in_theta = 1.741211 pi
 12'b110111101111: begin out_real=16'b0010110000001111; out_imag=16'b1101000110010101; end // in_theta = 1.741699 pi
 12'b110111110000: begin out_real=16'b0010110000100001; out_imag=16'b1101000110100110; end // in_theta = 1.742188 pi
 12'b110111110001: begin out_real=16'b0010110000110100; out_imag=16'b1101000110110111; end // in_theta = 1.742676 pi
 12'b110111110010: begin out_real=16'b0010110001000110; out_imag=16'b1101000111001001; end // in_theta = 1.743164 pi
 12'b110111110011: begin out_real=16'b0010110001011000; out_imag=16'b1101000111011010; end // in_theta = 1.743652 pi
 12'b110111110100: begin out_real=16'b0010110001101010; out_imag=16'b1101000111101011; end // in_theta = 1.744141 pi
 12'b110111110101: begin out_real=16'b0010110001111100; out_imag=16'b1101000111111101; end // in_theta = 1.744629 pi
 12'b110111110110: begin out_real=16'b0010110010001110; out_imag=16'b1101001000001110; end // in_theta = 1.745117 pi
 12'b110111110111: begin out_real=16'b0010110010100000; out_imag=16'b1101001000100000; end // in_theta = 1.745605 pi
 12'b110111111000: begin out_real=16'b0010110010110010; out_imag=16'b1101001000110001; end // in_theta = 1.746094 pi
 12'b110111111001: begin out_real=16'b0010110011000100; out_imag=16'b1101001001000011; end // in_theta = 1.746582 pi
 12'b110111111010: begin out_real=16'b0010110011010110; out_imag=16'b1101001001010101; end // in_theta = 1.747070 pi
 12'b110111111011: begin out_real=16'b0010110011101000; out_imag=16'b1101001001100110; end // in_theta = 1.747559 pi
 12'b110111111100: begin out_real=16'b0010110011111010; out_imag=16'b1101001001111000; end // in_theta = 1.748047 pi
 12'b110111111101: begin out_real=16'b0010110100001100; out_imag=16'b1101001010001010; end // in_theta = 1.748535 pi
 12'b110111111110: begin out_real=16'b0010110100011110; out_imag=16'b1101001010011011; end // in_theta = 1.749023 pi
 12'b110111111111: begin out_real=16'b0010110100101111; out_imag=16'b1101001010101101; end // in_theta = 1.749512 pi
 12'b111000000000: begin out_real=16'b0010110101000001; out_imag=16'b1101001010111111; end // in_theta = 1.750000 pi
 12'b111000000001: begin out_real=16'b0010110101010011; out_imag=16'b1101001011010001; end // in_theta = 1.750488 pi
 12'b111000000010: begin out_real=16'b0010110101100101; out_imag=16'b1101001011100010; end // in_theta = 1.750977 pi
 12'b111000000011: begin out_real=16'b0010110101110110; out_imag=16'b1101001011110100; end // in_theta = 1.751465 pi
 12'b111000000100: begin out_real=16'b0010110110001000; out_imag=16'b1101001100000110; end // in_theta = 1.751953 pi
 12'b111000000101: begin out_real=16'b0010110110011010; out_imag=16'b1101001100011000; end // in_theta = 1.752441 pi
 12'b111000000110: begin out_real=16'b0010110110101011; out_imag=16'b1101001100101010; end // in_theta = 1.752930 pi
 12'b111000000111: begin out_real=16'b0010110110111101; out_imag=16'b1101001100111100; end // in_theta = 1.753418 pi
 12'b111000001000: begin out_real=16'b0010110111001111; out_imag=16'b1101001101001110; end // in_theta = 1.753906 pi
 12'b111000001001: begin out_real=16'b0010110111100000; out_imag=16'b1101001101100000; end // in_theta = 1.754395 pi
 12'b111000001010: begin out_real=16'b0010110111110010; out_imag=16'b1101001101110010; end // in_theta = 1.754883 pi
 12'b111000001011: begin out_real=16'b0010111000000011; out_imag=16'b1101001110000100; end // in_theta = 1.755371 pi
 12'b111000001100: begin out_real=16'b0010111000010101; out_imag=16'b1101001110010110; end // in_theta = 1.755859 pi
 12'b111000001101: begin out_real=16'b0010111000100110; out_imag=16'b1101001110101000; end // in_theta = 1.756348 pi
 12'b111000001110: begin out_real=16'b0010111000110111; out_imag=16'b1101001110111010; end // in_theta = 1.756836 pi
 12'b111000001111: begin out_real=16'b0010111001001001; out_imag=16'b1101001111001100; end // in_theta = 1.757324 pi
 12'b111000010000: begin out_real=16'b0010111001011010; out_imag=16'b1101001111011111; end // in_theta = 1.757813 pi
 12'b111000010001: begin out_real=16'b0010111001101011; out_imag=16'b1101001111110001; end // in_theta = 1.758301 pi
 12'b111000010010: begin out_real=16'b0010111001111101; out_imag=16'b1101010000000011; end // in_theta = 1.758789 pi
 12'b111000010011: begin out_real=16'b0010111010001110; out_imag=16'b1101010000010101; end // in_theta = 1.759277 pi
 12'b111000010100: begin out_real=16'b0010111010011111; out_imag=16'b1101010000101000; end // in_theta = 1.759766 pi
 12'b111000010101: begin out_real=16'b0010111010110000; out_imag=16'b1101010000111010; end // in_theta = 1.760254 pi
 12'b111000010110: begin out_real=16'b0010111011000010; out_imag=16'b1101010001001100; end // in_theta = 1.760742 pi
 12'b111000010111: begin out_real=16'b0010111011010011; out_imag=16'b1101010001011111; end // in_theta = 1.761230 pi
 12'b111000011000: begin out_real=16'b0010111011100100; out_imag=16'b1101010001110001; end // in_theta = 1.761719 pi
 12'b111000011001: begin out_real=16'b0010111011110101; out_imag=16'b1101010010000011; end // in_theta = 1.762207 pi
 12'b111000011010: begin out_real=16'b0010111100000110; out_imag=16'b1101010010010110; end // in_theta = 1.762695 pi
 12'b111000011011: begin out_real=16'b0010111100010111; out_imag=16'b1101010010101000; end // in_theta = 1.763184 pi
 12'b111000011100: begin out_real=16'b0010111100101000; out_imag=16'b1101010010111011; end // in_theta = 1.763672 pi
 12'b111000011101: begin out_real=16'b0010111100111001; out_imag=16'b1101010011001101; end // in_theta = 1.764160 pi
 12'b111000011110: begin out_real=16'b0010111101001010; out_imag=16'b1101010011100000; end // in_theta = 1.764648 pi
 12'b111000011111: begin out_real=16'b0010111101011011; out_imag=16'b1101010011110011; end // in_theta = 1.765137 pi
 12'b111000100000: begin out_real=16'b0010111101101100; out_imag=16'b1101010100000101; end // in_theta = 1.765625 pi
 12'b111000100001: begin out_real=16'b0010111101111101; out_imag=16'b1101010100011000; end // in_theta = 1.766113 pi
 12'b111000100010: begin out_real=16'b0010111110001101; out_imag=16'b1101010100101010; end // in_theta = 1.766602 pi
 12'b111000100011: begin out_real=16'b0010111110011110; out_imag=16'b1101010100111101; end // in_theta = 1.767090 pi
 12'b111000100100: begin out_real=16'b0010111110101111; out_imag=16'b1101010101010000; end // in_theta = 1.767578 pi
 12'b111000100101: begin out_real=16'b0010111111000000; out_imag=16'b1101010101100011; end // in_theta = 1.768066 pi
 12'b111000100110: begin out_real=16'b0010111111010000; out_imag=16'b1101010101110101; end // in_theta = 1.768555 pi
 12'b111000100111: begin out_real=16'b0010111111100001; out_imag=16'b1101010110001000; end // in_theta = 1.769043 pi
 12'b111000101000: begin out_real=16'b0010111111110010; out_imag=16'b1101010110011011; end // in_theta = 1.769531 pi
 12'b111000101001: begin out_real=16'b0011000000000010; out_imag=16'b1101010110101110; end // in_theta = 1.770020 pi
 12'b111000101010: begin out_real=16'b0011000000010011; out_imag=16'b1101010111000001; end // in_theta = 1.770508 pi
 12'b111000101011: begin out_real=16'b0011000000100100; out_imag=16'b1101010111010100; end // in_theta = 1.770996 pi
 12'b111000101100: begin out_real=16'b0011000000110100; out_imag=16'b1101010111100110; end // in_theta = 1.771484 pi
 12'b111000101101: begin out_real=16'b0011000001000101; out_imag=16'b1101010111111001; end // in_theta = 1.771973 pi
 12'b111000101110: begin out_real=16'b0011000001010101; out_imag=16'b1101011000001100; end // in_theta = 1.772461 pi
 12'b111000101111: begin out_real=16'b0011000001100110; out_imag=16'b1101011000011111; end // in_theta = 1.772949 pi
 12'b111000110000: begin out_real=16'b0011000001110110; out_imag=16'b1101011000110010; end // in_theta = 1.773438 pi
 12'b111000110001: begin out_real=16'b0011000010000111; out_imag=16'b1101011001000101; end // in_theta = 1.773926 pi
 12'b111000110010: begin out_real=16'b0011000010010111; out_imag=16'b1101011001011001; end // in_theta = 1.774414 pi
 12'b111000110011: begin out_real=16'b0011000010100111; out_imag=16'b1101011001101100; end // in_theta = 1.774902 pi
 12'b111000110100: begin out_real=16'b0011000010111000; out_imag=16'b1101011001111111; end // in_theta = 1.775391 pi
 12'b111000110101: begin out_real=16'b0011000011001000; out_imag=16'b1101011010010010; end // in_theta = 1.775879 pi
 12'b111000110110: begin out_real=16'b0011000011011000; out_imag=16'b1101011010100101; end // in_theta = 1.776367 pi
 12'b111000110111: begin out_real=16'b0011000011101000; out_imag=16'b1101011010111000; end // in_theta = 1.776855 pi
 12'b111000111000: begin out_real=16'b0011000011111001; out_imag=16'b1101011011001011; end // in_theta = 1.777344 pi
 12'b111000111001: begin out_real=16'b0011000100001001; out_imag=16'b1101011011011111; end // in_theta = 1.777832 pi
 12'b111000111010: begin out_real=16'b0011000100011001; out_imag=16'b1101011011110010; end // in_theta = 1.778320 pi
 12'b111000111011: begin out_real=16'b0011000100101001; out_imag=16'b1101011100000101; end // in_theta = 1.778809 pi
 12'b111000111100: begin out_real=16'b0011000100111001; out_imag=16'b1101011100011001; end // in_theta = 1.779297 pi
 12'b111000111101: begin out_real=16'b0011000101001001; out_imag=16'b1101011100101100; end // in_theta = 1.779785 pi
 12'b111000111110: begin out_real=16'b0011000101011001; out_imag=16'b1101011100111111; end // in_theta = 1.780273 pi
 12'b111000111111: begin out_real=16'b0011000101101001; out_imag=16'b1101011101010011; end // in_theta = 1.780762 pi
 12'b111001000000: begin out_real=16'b0011000101111001; out_imag=16'b1101011101100110; end // in_theta = 1.781250 pi
 12'b111001000001: begin out_real=16'b0011000110001001; out_imag=16'b1101011101111010; end // in_theta = 1.781738 pi
 12'b111001000010: begin out_real=16'b0011000110011001; out_imag=16'b1101011110001101; end // in_theta = 1.782227 pi
 12'b111001000011: begin out_real=16'b0011000110101001; out_imag=16'b1101011110100000; end // in_theta = 1.782715 pi
 12'b111001000100: begin out_real=16'b0011000110111001; out_imag=16'b1101011110110100; end // in_theta = 1.783203 pi
 12'b111001000101: begin out_real=16'b0011000111001000; out_imag=16'b1101011111001000; end // in_theta = 1.783691 pi
 12'b111001000110: begin out_real=16'b0011000111011000; out_imag=16'b1101011111011011; end // in_theta = 1.784180 pi
 12'b111001000111: begin out_real=16'b0011000111101000; out_imag=16'b1101011111101111; end // in_theta = 1.784668 pi
 12'b111001001000: begin out_real=16'b0011000111111000; out_imag=16'b1101100000000010; end // in_theta = 1.785156 pi
 12'b111001001001: begin out_real=16'b0011001000000111; out_imag=16'b1101100000010110; end // in_theta = 1.785645 pi
 12'b111001001010: begin out_real=16'b0011001000010111; out_imag=16'b1101100000101010; end // in_theta = 1.786133 pi
 12'b111001001011: begin out_real=16'b0011001000100111; out_imag=16'b1101100000111101; end // in_theta = 1.786621 pi
 12'b111001001100: begin out_real=16'b0011001000110110; out_imag=16'b1101100001010001; end // in_theta = 1.787109 pi
 12'b111001001101: begin out_real=16'b0011001001000110; out_imag=16'b1101100001100101; end // in_theta = 1.787598 pi
 12'b111001001110: begin out_real=16'b0011001001010101; out_imag=16'b1101100001111000; end // in_theta = 1.788086 pi
 12'b111001001111: begin out_real=16'b0011001001100101; out_imag=16'b1101100010001100; end // in_theta = 1.788574 pi
 12'b111001010000: begin out_real=16'b0011001001110100; out_imag=16'b1101100010100000; end // in_theta = 1.789062 pi
 12'b111001010001: begin out_real=16'b0011001010000100; out_imag=16'b1101100010110100; end // in_theta = 1.789551 pi
 12'b111001010010: begin out_real=16'b0011001010010011; out_imag=16'b1101100011001000; end // in_theta = 1.790039 pi
 12'b111001010011: begin out_real=16'b0011001010100011; out_imag=16'b1101100011011100; end // in_theta = 1.790527 pi
 12'b111001010100: begin out_real=16'b0011001010110010; out_imag=16'b1101100011101111; end // in_theta = 1.791016 pi
 12'b111001010101: begin out_real=16'b0011001011000001; out_imag=16'b1101100100000011; end // in_theta = 1.791504 pi
 12'b111001010110: begin out_real=16'b0011001011010000; out_imag=16'b1101100100010111; end // in_theta = 1.791992 pi
 12'b111001010111: begin out_real=16'b0011001011100000; out_imag=16'b1101100100101011; end // in_theta = 1.792480 pi
 12'b111001011000: begin out_real=16'b0011001011101111; out_imag=16'b1101100100111111; end // in_theta = 1.792969 pi
 12'b111001011001: begin out_real=16'b0011001011111110; out_imag=16'b1101100101010011; end // in_theta = 1.793457 pi
 12'b111001011010: begin out_real=16'b0011001100001101; out_imag=16'b1101100101100111; end // in_theta = 1.793945 pi
 12'b111001011011: begin out_real=16'b0011001100011101; out_imag=16'b1101100101111011; end // in_theta = 1.794434 pi
 12'b111001011100: begin out_real=16'b0011001100101100; out_imag=16'b1101100110001111; end // in_theta = 1.794922 pi
 12'b111001011101: begin out_real=16'b0011001100111011; out_imag=16'b1101100110100100; end // in_theta = 1.795410 pi
 12'b111001011110: begin out_real=16'b0011001101001010; out_imag=16'b1101100110111000; end // in_theta = 1.795898 pi
 12'b111001011111: begin out_real=16'b0011001101011001; out_imag=16'b1101100111001100; end // in_theta = 1.796387 pi
 12'b111001100000: begin out_real=16'b0011001101101000; out_imag=16'b1101100111100000; end // in_theta = 1.796875 pi
 12'b111001100001: begin out_real=16'b0011001101110111; out_imag=16'b1101100111110100; end // in_theta = 1.797363 pi
 12'b111001100010: begin out_real=16'b0011001110000110; out_imag=16'b1101101000001000; end // in_theta = 1.797852 pi
 12'b111001100011: begin out_real=16'b0011001110010101; out_imag=16'b1101101000011101; end // in_theta = 1.798340 pi
 12'b111001100100: begin out_real=16'b0011001110100011; out_imag=16'b1101101000110001; end // in_theta = 1.798828 pi
 12'b111001100101: begin out_real=16'b0011001110110010; out_imag=16'b1101101001000101; end // in_theta = 1.799316 pi
 12'b111001100110: begin out_real=16'b0011001111000001; out_imag=16'b1101101001011010; end // in_theta = 1.799805 pi
 12'b111001100111: begin out_real=16'b0011001111010000; out_imag=16'b1101101001101110; end // in_theta = 1.800293 pi
 12'b111001101000: begin out_real=16'b0011001111011111; out_imag=16'b1101101010000010; end // in_theta = 1.800781 pi
 12'b111001101001: begin out_real=16'b0011001111101101; out_imag=16'b1101101010010111; end // in_theta = 1.801270 pi
 12'b111001101010: begin out_real=16'b0011001111111100; out_imag=16'b1101101010101011; end // in_theta = 1.801758 pi
 12'b111001101011: begin out_real=16'b0011010000001011; out_imag=16'b1101101010111111; end // in_theta = 1.802246 pi
 12'b111001101100: begin out_real=16'b0011010000011001; out_imag=16'b1101101011010100; end // in_theta = 1.802734 pi
 12'b111001101101: begin out_real=16'b0011010000101000; out_imag=16'b1101101011101000; end // in_theta = 1.803223 pi
 12'b111001101110: begin out_real=16'b0011010000110110; out_imag=16'b1101101011111101; end // in_theta = 1.803711 pi
 12'b111001101111: begin out_real=16'b0011010001000101; out_imag=16'b1101101100010001; end // in_theta = 1.804199 pi
 12'b111001110000: begin out_real=16'b0011010001010011; out_imag=16'b1101101100100110; end // in_theta = 1.804688 pi
 12'b111001110001: begin out_real=16'b0011010001100010; out_imag=16'b1101101100111011; end // in_theta = 1.805176 pi
 12'b111001110010: begin out_real=16'b0011010001110000; out_imag=16'b1101101101001111; end // in_theta = 1.805664 pi
 12'b111001110011: begin out_real=16'b0011010001111111; out_imag=16'b1101101101100100; end // in_theta = 1.806152 pi
 12'b111001110100: begin out_real=16'b0011010010001101; out_imag=16'b1101101101111000; end // in_theta = 1.806641 pi
 12'b111001110101: begin out_real=16'b0011010010011011; out_imag=16'b1101101110001101; end // in_theta = 1.807129 pi
 12'b111001110110: begin out_real=16'b0011010010101010; out_imag=16'b1101101110100010; end // in_theta = 1.807617 pi
 12'b111001110111: begin out_real=16'b0011010010111000; out_imag=16'b1101101110110110; end // in_theta = 1.808105 pi
 12'b111001111000: begin out_real=16'b0011010011000110; out_imag=16'b1101101111001011; end // in_theta = 1.808594 pi
 12'b111001111001: begin out_real=16'b0011010011010100; out_imag=16'b1101101111100000; end // in_theta = 1.809082 pi
 12'b111001111010: begin out_real=16'b0011010011100010; out_imag=16'b1101101111110101; end // in_theta = 1.809570 pi
 12'b111001111011: begin out_real=16'b0011010011110001; out_imag=16'b1101110000001001; end // in_theta = 1.810059 pi
 12'b111001111100: begin out_real=16'b0011010011111111; out_imag=16'b1101110000011110; end // in_theta = 1.810547 pi
 12'b111001111101: begin out_real=16'b0011010100001101; out_imag=16'b1101110000110011; end // in_theta = 1.811035 pi
 12'b111001111110: begin out_real=16'b0011010100011011; out_imag=16'b1101110001001000; end // in_theta = 1.811523 pi
 12'b111001111111: begin out_real=16'b0011010100101001; out_imag=16'b1101110001011101; end // in_theta = 1.812012 pi
 12'b111010000000: begin out_real=16'b0011010100110111; out_imag=16'b1101110001110010; end // in_theta = 1.812500 pi
 12'b111010000001: begin out_real=16'b0011010101000101; out_imag=16'b1101110010000110; end // in_theta = 1.812988 pi
 12'b111010000010: begin out_real=16'b0011010101010011; out_imag=16'b1101110010011011; end // in_theta = 1.813477 pi
 12'b111010000011: begin out_real=16'b0011010101100001; out_imag=16'b1101110010110000; end // in_theta = 1.813965 pi
 12'b111010000100: begin out_real=16'b0011010101101110; out_imag=16'b1101110011000101; end // in_theta = 1.814453 pi
 12'b111010000101: begin out_real=16'b0011010101111100; out_imag=16'b1101110011011010; end // in_theta = 1.814941 pi
 12'b111010000110: begin out_real=16'b0011010110001010; out_imag=16'b1101110011101111; end // in_theta = 1.815430 pi
 12'b111010000111: begin out_real=16'b0011010110011000; out_imag=16'b1101110100000100; end // in_theta = 1.815918 pi
 12'b111010001000: begin out_real=16'b0011010110100101; out_imag=16'b1101110100011001; end // in_theta = 1.816406 pi
 12'b111010001001: begin out_real=16'b0011010110110011; out_imag=16'b1101110100101110; end // in_theta = 1.816895 pi
 12'b111010001010: begin out_real=16'b0011010111000001; out_imag=16'b1101110101000100; end // in_theta = 1.817383 pi
 12'b111010001011: begin out_real=16'b0011010111001110; out_imag=16'b1101110101011001; end // in_theta = 1.817871 pi
 12'b111010001100: begin out_real=16'b0011010111011100; out_imag=16'b1101110101101110; end // in_theta = 1.818359 pi
 12'b111010001101: begin out_real=16'b0011010111101010; out_imag=16'b1101110110000011; end // in_theta = 1.818848 pi
 12'b111010001110: begin out_real=16'b0011010111110111; out_imag=16'b1101110110011000; end // in_theta = 1.819336 pi
 12'b111010001111: begin out_real=16'b0011011000000101; out_imag=16'b1101110110101101; end // in_theta = 1.819824 pi
 12'b111010010000: begin out_real=16'b0011011000010010; out_imag=16'b1101110111000011; end // in_theta = 1.820313 pi
 12'b111010010001: begin out_real=16'b0011011000100000; out_imag=16'b1101110111011000; end // in_theta = 1.820801 pi
 12'b111010010010: begin out_real=16'b0011011000101101; out_imag=16'b1101110111101101; end // in_theta = 1.821289 pi
 12'b111010010011: begin out_real=16'b0011011000111010; out_imag=16'b1101111000000010; end // in_theta = 1.821777 pi
 12'b111010010100: begin out_real=16'b0011011001001000; out_imag=16'b1101111000011000; end // in_theta = 1.822266 pi
 12'b111010010101: begin out_real=16'b0011011001010101; out_imag=16'b1101111000101101; end // in_theta = 1.822754 pi
 12'b111010010110: begin out_real=16'b0011011001100010; out_imag=16'b1101111001000010; end // in_theta = 1.823242 pi
 12'b111010010111: begin out_real=16'b0011011001101111; out_imag=16'b1101111001011000; end // in_theta = 1.823730 pi
 12'b111010011000: begin out_real=16'b0011011001111101; out_imag=16'b1101111001101101; end // in_theta = 1.824219 pi
 12'b111010011001: begin out_real=16'b0011011010001010; out_imag=16'b1101111010000011; end // in_theta = 1.824707 pi
 12'b111010011010: begin out_real=16'b0011011010010111; out_imag=16'b1101111010011000; end // in_theta = 1.825195 pi
 12'b111010011011: begin out_real=16'b0011011010100100; out_imag=16'b1101111010101101; end // in_theta = 1.825684 pi
 12'b111010011100: begin out_real=16'b0011011010110001; out_imag=16'b1101111011000011; end // in_theta = 1.826172 pi
 12'b111010011101: begin out_real=16'b0011011010111110; out_imag=16'b1101111011011000; end // in_theta = 1.826660 pi
 12'b111010011110: begin out_real=16'b0011011011001011; out_imag=16'b1101111011101110; end // in_theta = 1.827148 pi
 12'b111010011111: begin out_real=16'b0011011011011000; out_imag=16'b1101111100000011; end // in_theta = 1.827637 pi
 12'b111010100000: begin out_real=16'b0011011011100101; out_imag=16'b1101111100011001; end // in_theta = 1.828125 pi
 12'b111010100001: begin out_real=16'b0011011011110010; out_imag=16'b1101111100101111; end // in_theta = 1.828613 pi
 12'b111010100010: begin out_real=16'b0011011011111111; out_imag=16'b1101111101000100; end // in_theta = 1.829102 pi
 12'b111010100011: begin out_real=16'b0011011100001100; out_imag=16'b1101111101011010; end // in_theta = 1.829590 pi
 12'b111010100100: begin out_real=16'b0011011100011000; out_imag=16'b1101111101101111; end // in_theta = 1.830078 pi
 12'b111010100101: begin out_real=16'b0011011100100101; out_imag=16'b1101111110000101; end // in_theta = 1.830566 pi
 12'b111010100110: begin out_real=16'b0011011100110010; out_imag=16'b1101111110011011; end // in_theta = 1.831055 pi
 12'b111010100111: begin out_real=16'b0011011100111111; out_imag=16'b1101111110110000; end // in_theta = 1.831543 pi
 12'b111010101000: begin out_real=16'b0011011101001011; out_imag=16'b1101111111000110; end // in_theta = 1.832031 pi
 12'b111010101001: begin out_real=16'b0011011101011000; out_imag=16'b1101111111011100; end // in_theta = 1.832520 pi
 12'b111010101010: begin out_real=16'b0011011101100101; out_imag=16'b1101111111110001; end // in_theta = 1.833008 pi
 12'b111010101011: begin out_real=16'b0011011101110001; out_imag=16'b1110000000000111; end // in_theta = 1.833496 pi
 12'b111010101100: begin out_real=16'b0011011101111110; out_imag=16'b1110000000011101; end // in_theta = 1.833984 pi
 12'b111010101101: begin out_real=16'b0011011110001010; out_imag=16'b1110000000110011; end // in_theta = 1.834473 pi
 12'b111010101110: begin out_real=16'b0011011110010111; out_imag=16'b1110000001001001; end // in_theta = 1.834961 pi
 12'b111010101111: begin out_real=16'b0011011110100011; out_imag=16'b1110000001011110; end // in_theta = 1.835449 pi
 12'b111010110000: begin out_real=16'b0011011110110000; out_imag=16'b1110000001110100; end // in_theta = 1.835938 pi
 12'b111010110001: begin out_real=16'b0011011110111100; out_imag=16'b1110000010001010; end // in_theta = 1.836426 pi
 12'b111010110010: begin out_real=16'b0011011111001000; out_imag=16'b1110000010100000; end // in_theta = 1.836914 pi
 12'b111010110011: begin out_real=16'b0011011111010101; out_imag=16'b1110000010110110; end // in_theta = 1.837402 pi
 12'b111010110100: begin out_real=16'b0011011111100001; out_imag=16'b1110000011001100; end // in_theta = 1.837891 pi
 12'b111010110101: begin out_real=16'b0011011111101101; out_imag=16'b1110000011100010; end // in_theta = 1.838379 pi
 12'b111010110110: begin out_real=16'b0011011111111001; out_imag=16'b1110000011111000; end // in_theta = 1.838867 pi
 12'b111010110111: begin out_real=16'b0011100000000101; out_imag=16'b1110000100001110; end // in_theta = 1.839355 pi
 12'b111010111000: begin out_real=16'b0011100000010010; out_imag=16'b1110000100100100; end // in_theta = 1.839844 pi
 12'b111010111001: begin out_real=16'b0011100000011110; out_imag=16'b1110000100111010; end // in_theta = 1.840332 pi
 12'b111010111010: begin out_real=16'b0011100000101010; out_imag=16'b1110000101010000; end // in_theta = 1.840820 pi
 12'b111010111011: begin out_real=16'b0011100000110110; out_imag=16'b1110000101100110; end // in_theta = 1.841309 pi
 12'b111010111100: begin out_real=16'b0011100001000010; out_imag=16'b1110000101111100; end // in_theta = 1.841797 pi
 12'b111010111101: begin out_real=16'b0011100001001110; out_imag=16'b1110000110010010; end // in_theta = 1.842285 pi
 12'b111010111110: begin out_real=16'b0011100001011010; out_imag=16'b1110000110101000; end // in_theta = 1.842773 pi
 12'b111010111111: begin out_real=16'b0011100001100110; out_imag=16'b1110000110111110; end // in_theta = 1.843262 pi
 12'b111011000000: begin out_real=16'b0011100001110001; out_imag=16'b1110000111010101; end // in_theta = 1.843750 pi
 12'b111011000001: begin out_real=16'b0011100001111101; out_imag=16'b1110000111101011; end // in_theta = 1.844238 pi
 12'b111011000010: begin out_real=16'b0011100010001001; out_imag=16'b1110001000000001; end // in_theta = 1.844727 pi
 12'b111011000011: begin out_real=16'b0011100010010101; out_imag=16'b1110001000010111; end // in_theta = 1.845215 pi
 12'b111011000100: begin out_real=16'b0011100010100001; out_imag=16'b1110001000101101; end // in_theta = 1.845703 pi
 12'b111011000101: begin out_real=16'b0011100010101100; out_imag=16'b1110001001000100; end // in_theta = 1.846191 pi
 12'b111011000110: begin out_real=16'b0011100010111000; out_imag=16'b1110001001011010; end // in_theta = 1.846680 pi
 12'b111011000111: begin out_real=16'b0011100011000011; out_imag=16'b1110001001110000; end // in_theta = 1.847168 pi
 12'b111011001000: begin out_real=16'b0011100011001111; out_imag=16'b1110001010000111; end // in_theta = 1.847656 pi
 12'b111011001001: begin out_real=16'b0011100011011011; out_imag=16'b1110001010011101; end // in_theta = 1.848145 pi
 12'b111011001010: begin out_real=16'b0011100011100110; out_imag=16'b1110001010110011; end // in_theta = 1.848633 pi
 12'b111011001011: begin out_real=16'b0011100011110010; out_imag=16'b1110001011001010; end // in_theta = 1.849121 pi
 12'b111011001100: begin out_real=16'b0011100011111101; out_imag=16'b1110001011100000; end // in_theta = 1.849609 pi
 12'b111011001101: begin out_real=16'b0011100100001001; out_imag=16'b1110001011110110; end // in_theta = 1.850098 pi
 12'b111011001110: begin out_real=16'b0011100100010100; out_imag=16'b1110001100001101; end // in_theta = 1.850586 pi
 12'b111011001111: begin out_real=16'b0011100100011111; out_imag=16'b1110001100100011; end // in_theta = 1.851074 pi
 12'b111011010000: begin out_real=16'b0011100100101011; out_imag=16'b1110001100111010; end // in_theta = 1.851563 pi
 12'b111011010001: begin out_real=16'b0011100100110110; out_imag=16'b1110001101010000; end // in_theta = 1.852051 pi
 12'b111011010010: begin out_real=16'b0011100101000001; out_imag=16'b1110001101100111; end // in_theta = 1.852539 pi
 12'b111011010011: begin out_real=16'b0011100101001100; out_imag=16'b1110001101111101; end // in_theta = 1.853027 pi
 12'b111011010100: begin out_real=16'b0011100101011000; out_imag=16'b1110001110010100; end // in_theta = 1.853516 pi
 12'b111011010101: begin out_real=16'b0011100101100011; out_imag=16'b1110001110101010; end // in_theta = 1.854004 pi
 12'b111011010110: begin out_real=16'b0011100101101110; out_imag=16'b1110001111000001; end // in_theta = 1.854492 pi
 12'b111011010111: begin out_real=16'b0011100101111001; out_imag=16'b1110001111010111; end // in_theta = 1.854980 pi
 12'b111011011000: begin out_real=16'b0011100110000100; out_imag=16'b1110001111101110; end // in_theta = 1.855469 pi
 12'b111011011001: begin out_real=16'b0011100110001111; out_imag=16'b1110010000000100; end // in_theta = 1.855957 pi
 12'b111011011010: begin out_real=16'b0011100110011010; out_imag=16'b1110010000011011; end // in_theta = 1.856445 pi
 12'b111011011011: begin out_real=16'b0011100110100101; out_imag=16'b1110010000110010; end // in_theta = 1.856934 pi
 12'b111011011100: begin out_real=16'b0011100110110000; out_imag=16'b1110010001001000; end // in_theta = 1.857422 pi
 12'b111011011101: begin out_real=16'b0011100110111011; out_imag=16'b1110010001011111; end // in_theta = 1.857910 pi
 12'b111011011110: begin out_real=16'b0011100111000101; out_imag=16'b1110010001110110; end // in_theta = 1.858398 pi
 12'b111011011111: begin out_real=16'b0011100111010000; out_imag=16'b1110010010001100; end // in_theta = 1.858887 pi
 12'b111011100000: begin out_real=16'b0011100111011011; out_imag=16'b1110010010100011; end // in_theta = 1.859375 pi
 12'b111011100001: begin out_real=16'b0011100111100110; out_imag=16'b1110010010111010; end // in_theta = 1.859863 pi
 12'b111011100010: begin out_real=16'b0011100111110000; out_imag=16'b1110010011010000; end // in_theta = 1.860352 pi
 12'b111011100011: begin out_real=16'b0011100111111011; out_imag=16'b1110010011100111; end // in_theta = 1.860840 pi
 12'b111011100100: begin out_real=16'b0011101000000110; out_imag=16'b1110010011111110; end // in_theta = 1.861328 pi
 12'b111011100101: begin out_real=16'b0011101000010000; out_imag=16'b1110010100010101; end // in_theta = 1.861816 pi
 12'b111011100110: begin out_real=16'b0011101000011011; out_imag=16'b1110010100101100; end // in_theta = 1.862305 pi
 12'b111011100111: begin out_real=16'b0011101000100101; out_imag=16'b1110010101000010; end // in_theta = 1.862793 pi
 12'b111011101000: begin out_real=16'b0011101000110000; out_imag=16'b1110010101011001; end // in_theta = 1.863281 pi
 12'b111011101001: begin out_real=16'b0011101000111010; out_imag=16'b1110010101110000; end // in_theta = 1.863770 pi
 12'b111011101010: begin out_real=16'b0011101001000101; out_imag=16'b1110010110000111; end // in_theta = 1.864258 pi
 12'b111011101011: begin out_real=16'b0011101001001111; out_imag=16'b1110010110011110; end // in_theta = 1.864746 pi
 12'b111011101100: begin out_real=16'b0011101001011001; out_imag=16'b1110010110110101; end // in_theta = 1.865234 pi
 12'b111011101101: begin out_real=16'b0011101001100100; out_imag=16'b1110010111001100; end // in_theta = 1.865723 pi
 12'b111011101110: begin out_real=16'b0011101001101110; out_imag=16'b1110010111100011; end // in_theta = 1.866211 pi
 12'b111011101111: begin out_real=16'b0011101001111000; out_imag=16'b1110010111111010; end // in_theta = 1.866699 pi
 12'b111011110000: begin out_real=16'b0011101010000010; out_imag=16'b1110011000010001; end // in_theta = 1.867187 pi
 12'b111011110001: begin out_real=16'b0011101010001101; out_imag=16'b1110011000101000; end // in_theta = 1.867676 pi
 12'b111011110010: begin out_real=16'b0011101010010111; out_imag=16'b1110011000111111; end // in_theta = 1.868164 pi
 12'b111011110011: begin out_real=16'b0011101010100001; out_imag=16'b1110011001010110; end // in_theta = 1.868652 pi
 12'b111011110100: begin out_real=16'b0011101010101011; out_imag=16'b1110011001101101; end // in_theta = 1.869141 pi
 12'b111011110101: begin out_real=16'b0011101010110101; out_imag=16'b1110011010000100; end // in_theta = 1.869629 pi
 12'b111011110110: begin out_real=16'b0011101010111111; out_imag=16'b1110011010011011; end // in_theta = 1.870117 pi
 12'b111011110111: begin out_real=16'b0011101011001001; out_imag=16'b1110011010110010; end // in_theta = 1.870605 pi
 12'b111011111000: begin out_real=16'b0011101011010011; out_imag=16'b1110011011001001; end // in_theta = 1.871094 pi
 12'b111011111001: begin out_real=16'b0011101011011101; out_imag=16'b1110011011100000; end // in_theta = 1.871582 pi
 12'b111011111010: begin out_real=16'b0011101011100110; out_imag=16'b1110011011110111; end // in_theta = 1.872070 pi
 12'b111011111011: begin out_real=16'b0011101011110000; out_imag=16'b1110011100001110; end // in_theta = 1.872559 pi
 12'b111011111100: begin out_real=16'b0011101011111010; out_imag=16'b1110011100100101; end // in_theta = 1.873047 pi
 12'b111011111101: begin out_real=16'b0011101100000100; out_imag=16'b1110011100111101; end // in_theta = 1.873535 pi
 12'b111011111110: begin out_real=16'b0011101100001110; out_imag=16'b1110011101010100; end // in_theta = 1.874023 pi
 12'b111011111111: begin out_real=16'b0011101100010111; out_imag=16'b1110011101101011; end // in_theta = 1.874512 pi
 12'b111100000000: begin out_real=16'b0011101100100001; out_imag=16'b1110011110000010; end // in_theta = 1.875000 pi
 12'b111100000001: begin out_real=16'b0011101100101010; out_imag=16'b1110011110011001; end // in_theta = 1.875488 pi
 12'b111100000010: begin out_real=16'b0011101100110100; out_imag=16'b1110011110110001; end // in_theta = 1.875977 pi
 12'b111100000011: begin out_real=16'b0011101100111110; out_imag=16'b1110011111001000; end // in_theta = 1.876465 pi
 12'b111100000100: begin out_real=16'b0011101101000111; out_imag=16'b1110011111011111; end // in_theta = 1.876953 pi
 12'b111100000101: begin out_real=16'b0011101101010000; out_imag=16'b1110011111110110; end // in_theta = 1.877441 pi
 12'b111100000110: begin out_real=16'b0011101101011010; out_imag=16'b1110100000001110; end // in_theta = 1.877930 pi
 12'b111100000111: begin out_real=16'b0011101101100011; out_imag=16'b1110100000100101; end // in_theta = 1.878418 pi
 12'b111100001000: begin out_real=16'b0011101101101101; out_imag=16'b1110100000111100; end // in_theta = 1.878906 pi
 12'b111100001001: begin out_real=16'b0011101101110110; out_imag=16'b1110100001010100; end // in_theta = 1.879395 pi
 12'b111100001010: begin out_real=16'b0011101101111111; out_imag=16'b1110100001101011; end // in_theta = 1.879883 pi
 12'b111100001011: begin out_real=16'b0011101110001000; out_imag=16'b1110100010000010; end // in_theta = 1.880371 pi
 12'b111100001100: begin out_real=16'b0011101110010010; out_imag=16'b1110100010011010; end // in_theta = 1.880859 pi
 12'b111100001101: begin out_real=16'b0011101110011011; out_imag=16'b1110100010110001; end // in_theta = 1.881348 pi
 12'b111100001110: begin out_real=16'b0011101110100100; out_imag=16'b1110100011001001; end // in_theta = 1.881836 pi
 12'b111100001111: begin out_real=16'b0011101110101101; out_imag=16'b1110100011100000; end // in_theta = 1.882324 pi
 12'b111100010000: begin out_real=16'b0011101110110110; out_imag=16'b1110100011110111; end // in_theta = 1.882813 pi
 12'b111100010001: begin out_real=16'b0011101110111111; out_imag=16'b1110100100001111; end // in_theta = 1.883301 pi
 12'b111100010010: begin out_real=16'b0011101111001000; out_imag=16'b1110100100100110; end // in_theta = 1.883789 pi
 12'b111100010011: begin out_real=16'b0011101111010001; out_imag=16'b1110100100111110; end // in_theta = 1.884277 pi
 12'b111100010100: begin out_real=16'b0011101111011010; out_imag=16'b1110100101010101; end // in_theta = 1.884766 pi
 12'b111100010101: begin out_real=16'b0011101111100011; out_imag=16'b1110100101101101; end // in_theta = 1.885254 pi
 12'b111100010110: begin out_real=16'b0011101111101100; out_imag=16'b1110100110000100; end // in_theta = 1.885742 pi
 12'b111100010111: begin out_real=16'b0011101111110101; out_imag=16'b1110100110011100; end // in_theta = 1.886230 pi
 12'b111100011000: begin out_real=16'b0011101111111101; out_imag=16'b1110100110110100; end // in_theta = 1.886719 pi
 12'b111100011001: begin out_real=16'b0011110000000110; out_imag=16'b1110100111001011; end // in_theta = 1.887207 pi
 12'b111100011010: begin out_real=16'b0011110000001111; out_imag=16'b1110100111100011; end // in_theta = 1.887695 pi
 12'b111100011011: begin out_real=16'b0011110000010111; out_imag=16'b1110100111111010; end // in_theta = 1.888184 pi
 12'b111100011100: begin out_real=16'b0011110000100000; out_imag=16'b1110101000010010; end // in_theta = 1.888672 pi
 12'b111100011101: begin out_real=16'b0011110000101001; out_imag=16'b1110101000101001; end // in_theta = 1.889160 pi
 12'b111100011110: begin out_real=16'b0011110000110001; out_imag=16'b1110101001000001; end // in_theta = 1.889648 pi
 12'b111100011111: begin out_real=16'b0011110000111010; out_imag=16'b1110101001011001; end // in_theta = 1.890137 pi
 12'b111100100000: begin out_real=16'b0011110001000010; out_imag=16'b1110101001110000; end // in_theta = 1.890625 pi
 12'b111100100001: begin out_real=16'b0011110001001011; out_imag=16'b1110101010001000; end // in_theta = 1.891113 pi
 12'b111100100010: begin out_real=16'b0011110001010011; out_imag=16'b1110101010100000; end // in_theta = 1.891602 pi
 12'b111100100011: begin out_real=16'b0011110001011011; out_imag=16'b1110101010110111; end // in_theta = 1.892090 pi
 12'b111100100100: begin out_real=16'b0011110001100100; out_imag=16'b1110101011001111; end // in_theta = 1.892578 pi
 12'b111100100101: begin out_real=16'b0011110001101100; out_imag=16'b1110101011100111; end // in_theta = 1.893066 pi
 12'b111100100110: begin out_real=16'b0011110001110100; out_imag=16'b1110101011111111; end // in_theta = 1.893555 pi
 12'b111100100111: begin out_real=16'b0011110001111101; out_imag=16'b1110101100010110; end // in_theta = 1.894043 pi
 12'b111100101000: begin out_real=16'b0011110010000101; out_imag=16'b1110101100101110; end // in_theta = 1.894531 pi
 12'b111100101001: begin out_real=16'b0011110010001101; out_imag=16'b1110101101000110; end // in_theta = 1.895020 pi
 12'b111100101010: begin out_real=16'b0011110010010101; out_imag=16'b1110101101011110; end // in_theta = 1.895508 pi
 12'b111100101011: begin out_real=16'b0011110010011101; out_imag=16'b1110101101110101; end // in_theta = 1.895996 pi
 12'b111100101100: begin out_real=16'b0011110010100101; out_imag=16'b1110101110001101; end // in_theta = 1.896484 pi
 12'b111100101101: begin out_real=16'b0011110010101101; out_imag=16'b1110101110100101; end // in_theta = 1.896973 pi
 12'b111100101110: begin out_real=16'b0011110010110101; out_imag=16'b1110101110111101; end // in_theta = 1.897461 pi
 12'b111100101111: begin out_real=16'b0011110010111101; out_imag=16'b1110101111010101; end // in_theta = 1.897949 pi
 12'b111100110000: begin out_real=16'b0011110011000101; out_imag=16'b1110101111101101; end // in_theta = 1.898438 pi
 12'b111100110001: begin out_real=16'b0011110011001101; out_imag=16'b1110110000000101; end // in_theta = 1.898926 pi
 12'b111100110010: begin out_real=16'b0011110011010101; out_imag=16'b1110110000011100; end // in_theta = 1.899414 pi
 12'b111100110011: begin out_real=16'b0011110011011101; out_imag=16'b1110110000110100; end // in_theta = 1.899902 pi
 12'b111100110100: begin out_real=16'b0011110011100100; out_imag=16'b1110110001001100; end // in_theta = 1.900391 pi
 12'b111100110101: begin out_real=16'b0011110011101100; out_imag=16'b1110110001100100; end // in_theta = 1.900879 pi
 12'b111100110110: begin out_real=16'b0011110011110100; out_imag=16'b1110110001111100; end // in_theta = 1.901367 pi
 12'b111100110111: begin out_real=16'b0011110011111011; out_imag=16'b1110110010010100; end // in_theta = 1.901855 pi
 12'b111100111000: begin out_real=16'b0011110100000011; out_imag=16'b1110110010101100; end // in_theta = 1.902344 pi
 12'b111100111001: begin out_real=16'b0011110100001011; out_imag=16'b1110110011000100; end // in_theta = 1.902832 pi
 12'b111100111010: begin out_real=16'b0011110100010010; out_imag=16'b1110110011011100; end // in_theta = 1.903320 pi
 12'b111100111011: begin out_real=16'b0011110100011010; out_imag=16'b1110110011110100; end // in_theta = 1.903809 pi
 12'b111100111100: begin out_real=16'b0011110100100001; out_imag=16'b1110110100001100; end // in_theta = 1.904297 pi
 12'b111100111101: begin out_real=16'b0011110100101000; out_imag=16'b1110110100100100; end // in_theta = 1.904785 pi
 12'b111100111110: begin out_real=16'b0011110100110000; out_imag=16'b1110110100111100; end // in_theta = 1.905273 pi
 12'b111100111111: begin out_real=16'b0011110100110111; out_imag=16'b1110110101010100; end // in_theta = 1.905762 pi
 12'b111101000000: begin out_real=16'b0011110100111111; out_imag=16'b1110110101101100; end // in_theta = 1.906250 pi
 12'b111101000001: begin out_real=16'b0011110101000110; out_imag=16'b1110110110000100; end // in_theta = 1.906738 pi
 12'b111101000010: begin out_real=16'b0011110101001101; out_imag=16'b1110110110011100; end // in_theta = 1.907227 pi
 12'b111101000011: begin out_real=16'b0011110101010100; out_imag=16'b1110110110110100; end // in_theta = 1.907715 pi
 12'b111101000100: begin out_real=16'b0011110101011011; out_imag=16'b1110110111001100; end // in_theta = 1.908203 pi
 12'b111101000101: begin out_real=16'b0011110101100011; out_imag=16'b1110110111100100; end // in_theta = 1.908691 pi
 12'b111101000110: begin out_real=16'b0011110101101010; out_imag=16'b1110110111111100; end // in_theta = 1.909180 pi
 12'b111101000111: begin out_real=16'b0011110101110001; out_imag=16'b1110111000010101; end // in_theta = 1.909668 pi
 12'b111101001000: begin out_real=16'b0011110101111000; out_imag=16'b1110111000101101; end // in_theta = 1.910156 pi
 12'b111101001001: begin out_real=16'b0011110101111111; out_imag=16'b1110111001000101; end // in_theta = 1.910645 pi
 12'b111101001010: begin out_real=16'b0011110110000110; out_imag=16'b1110111001011101; end // in_theta = 1.911133 pi
 12'b111101001011: begin out_real=16'b0011110110001101; out_imag=16'b1110111001110101; end // in_theta = 1.911621 pi
 12'b111101001100: begin out_real=16'b0011110110010011; out_imag=16'b1110111010001101; end // in_theta = 1.912109 pi
 12'b111101001101: begin out_real=16'b0011110110011010; out_imag=16'b1110111010100110; end // in_theta = 1.912598 pi
 12'b111101001110: begin out_real=16'b0011110110100001; out_imag=16'b1110111010111110; end // in_theta = 1.913086 pi
 12'b111101001111: begin out_real=16'b0011110110101000; out_imag=16'b1110111011010110; end // in_theta = 1.913574 pi
 12'b111101010000: begin out_real=16'b0011110110101111; out_imag=16'b1110111011101110; end // in_theta = 1.914063 pi
 12'b111101010001: begin out_real=16'b0011110110110101; out_imag=16'b1110111100000110; end // in_theta = 1.914551 pi
 12'b111101010010: begin out_real=16'b0011110110111100; out_imag=16'b1110111100011111; end // in_theta = 1.915039 pi
 12'b111101010011: begin out_real=16'b0011110111000010; out_imag=16'b1110111100110111; end // in_theta = 1.915527 pi
 12'b111101010100: begin out_real=16'b0011110111001001; out_imag=16'b1110111101001111; end // in_theta = 1.916016 pi
 12'b111101010101: begin out_real=16'b0011110111010000; out_imag=16'b1110111101100111; end // in_theta = 1.916504 pi
 12'b111101010110: begin out_real=16'b0011110111010110; out_imag=16'b1110111110000000; end // in_theta = 1.916992 pi
 12'b111101010111: begin out_real=16'b0011110111011101; out_imag=16'b1110111110011000; end // in_theta = 1.917480 pi
 12'b111101011000: begin out_real=16'b0011110111100011; out_imag=16'b1110111110110000; end // in_theta = 1.917969 pi
 12'b111101011001: begin out_real=16'b0011110111101001; out_imag=16'b1110111111001001; end // in_theta = 1.918457 pi
 12'b111101011010: begin out_real=16'b0011110111110000; out_imag=16'b1110111111100001; end // in_theta = 1.918945 pi
 12'b111101011011: begin out_real=16'b0011110111110110; out_imag=16'b1110111111111001; end // in_theta = 1.919434 pi
 12'b111101011100: begin out_real=16'b0011110111111100; out_imag=16'b1111000000010010; end // in_theta = 1.919922 pi
 12'b111101011101: begin out_real=16'b0011111000000011; out_imag=16'b1111000000101010; end // in_theta = 1.920410 pi
 12'b111101011110: begin out_real=16'b0011111000001001; out_imag=16'b1111000001000010; end // in_theta = 1.920898 pi
 12'b111101011111: begin out_real=16'b0011111000001111; out_imag=16'b1111000001011011; end // in_theta = 1.921387 pi
 12'b111101100000: begin out_real=16'b0011111000010101; out_imag=16'b1111000001110011; end // in_theta = 1.921875 pi
 12'b111101100001: begin out_real=16'b0011111000011011; out_imag=16'b1111000010001011; end // in_theta = 1.922363 pi
 12'b111101100010: begin out_real=16'b0011111000100001; out_imag=16'b1111000010100100; end // in_theta = 1.922852 pi
 12'b111101100011: begin out_real=16'b0011111000100111; out_imag=16'b1111000010111100; end // in_theta = 1.923340 pi
 12'b111101100100: begin out_real=16'b0011111000101101; out_imag=16'b1111000011010101; end // in_theta = 1.923828 pi
 12'b111101100101: begin out_real=16'b0011111000110011; out_imag=16'b1111000011101101; end // in_theta = 1.924316 pi
 12'b111101100110: begin out_real=16'b0011111000111001; out_imag=16'b1111000100000101; end // in_theta = 1.924805 pi
 12'b111101100111: begin out_real=16'b0011111000111111; out_imag=16'b1111000100011110; end // in_theta = 1.925293 pi
 12'b111101101000: begin out_real=16'b0011111001000101; out_imag=16'b1111000100110110; end // in_theta = 1.925781 pi
 12'b111101101001: begin out_real=16'b0011111001001010; out_imag=16'b1111000101001111; end // in_theta = 1.926270 pi
 12'b111101101010: begin out_real=16'b0011111001010000; out_imag=16'b1111000101100111; end // in_theta = 1.926758 pi
 12'b111101101011: begin out_real=16'b0011111001010110; out_imag=16'b1111000110000000; end // in_theta = 1.927246 pi
 12'b111101101100: begin out_real=16'b0011111001011100; out_imag=16'b1111000110011000; end // in_theta = 1.927734 pi
 12'b111101101101: begin out_real=16'b0011111001100001; out_imag=16'b1111000110110001; end // in_theta = 1.928223 pi
 12'b111101101110: begin out_real=16'b0011111001100111; out_imag=16'b1111000111001001; end // in_theta = 1.928711 pi
 12'b111101101111: begin out_real=16'b0011111001101100; out_imag=16'b1111000111100010; end // in_theta = 1.929199 pi
 12'b111101110000: begin out_real=16'b0011111001110010; out_imag=16'b1111000111111010; end // in_theta = 1.929688 pi
 12'b111101110001: begin out_real=16'b0011111001110111; out_imag=16'b1111001000010011; end // in_theta = 1.930176 pi
 12'b111101110010: begin out_real=16'b0011111001111101; out_imag=16'b1111001000101011; end // in_theta = 1.930664 pi
 12'b111101110011: begin out_real=16'b0011111010000010; out_imag=16'b1111001001000100; end // in_theta = 1.931152 pi
 12'b111101110100: begin out_real=16'b0011111010001000; out_imag=16'b1111001001011100; end // in_theta = 1.931641 pi
 12'b111101110101: begin out_real=16'b0011111010001101; out_imag=16'b1111001001110101; end // in_theta = 1.932129 pi
 12'b111101110110: begin out_real=16'b0011111010010010; out_imag=16'b1111001010001110; end // in_theta = 1.932617 pi
 12'b111101110111: begin out_real=16'b0011111010011000; out_imag=16'b1111001010100110; end // in_theta = 1.933105 pi
 12'b111101111000: begin out_real=16'b0011111010011101; out_imag=16'b1111001010111111; end // in_theta = 1.933594 pi
 12'b111101111001: begin out_real=16'b0011111010100010; out_imag=16'b1111001011010111; end // in_theta = 1.934082 pi
 12'b111101111010: begin out_real=16'b0011111010100111; out_imag=16'b1111001011110000; end // in_theta = 1.934570 pi
 12'b111101111011: begin out_real=16'b0011111010101100; out_imag=16'b1111001100001000; end // in_theta = 1.935059 pi
 12'b111101111100: begin out_real=16'b0011111010110001; out_imag=16'b1111001100100001; end // in_theta = 1.935547 pi
 12'b111101111101: begin out_real=16'b0011111010110110; out_imag=16'b1111001100111010; end // in_theta = 1.936035 pi
 12'b111101111110: begin out_real=16'b0011111010111011; out_imag=16'b1111001101010010; end // in_theta = 1.936523 pi
 12'b111101111111: begin out_real=16'b0011111011000000; out_imag=16'b1111001101101011; end // in_theta = 1.937012 pi
 12'b111110000000: begin out_real=16'b0011111011000101; out_imag=16'b1111001110000100; end // in_theta = 1.937500 pi
 12'b111110000001: begin out_real=16'b0011111011001010; out_imag=16'b1111001110011100; end // in_theta = 1.937988 pi
 12'b111110000010: begin out_real=16'b0011111011001111; out_imag=16'b1111001110110101; end // in_theta = 1.938477 pi
 12'b111110000011: begin out_real=16'b0011111011010100; out_imag=16'b1111001111001110; end // in_theta = 1.938965 pi
 12'b111110000100: begin out_real=16'b0011111011011000; out_imag=16'b1111001111100110; end // in_theta = 1.939453 pi
 12'b111110000101: begin out_real=16'b0011111011011101; out_imag=16'b1111001111111111; end // in_theta = 1.939941 pi
 12'b111110000110: begin out_real=16'b0011111011100010; out_imag=16'b1111010000011000; end // in_theta = 1.940430 pi
 12'b111110000111: begin out_real=16'b0011111011100111; out_imag=16'b1111010000110000; end // in_theta = 1.940918 pi
 12'b111110001000: begin out_real=16'b0011111011101011; out_imag=16'b1111010001001001; end // in_theta = 1.941406 pi
 12'b111110001001: begin out_real=16'b0011111011110000; out_imag=16'b1111010001100010; end // in_theta = 1.941895 pi
 12'b111110001010: begin out_real=16'b0011111011110100; out_imag=16'b1111010001111011; end // in_theta = 1.942383 pi
 12'b111110001011: begin out_real=16'b0011111011111001; out_imag=16'b1111010010010011; end // in_theta = 1.942871 pi
 12'b111110001100: begin out_real=16'b0011111011111101; out_imag=16'b1111010010101100; end // in_theta = 1.943359 pi
 12'b111110001101: begin out_real=16'b0011111100000010; out_imag=16'b1111010011000101; end // in_theta = 1.943848 pi
 12'b111110001110: begin out_real=16'b0011111100000110; out_imag=16'b1111010011011101; end // in_theta = 1.944336 pi
 12'b111110001111: begin out_real=16'b0011111100001010; out_imag=16'b1111010011110110; end // in_theta = 1.944824 pi
 12'b111110010000: begin out_real=16'b0011111100001111; out_imag=16'b1111010100001111; end // in_theta = 1.945313 pi
 12'b111110010001: begin out_real=16'b0011111100010011; out_imag=16'b1111010100101000; end // in_theta = 1.945801 pi
 12'b111110010010: begin out_real=16'b0011111100010111; out_imag=16'b1111010101000000; end // in_theta = 1.946289 pi
 12'b111110010011: begin out_real=16'b0011111100011100; out_imag=16'b1111010101011001; end // in_theta = 1.946777 pi
 12'b111110010100: begin out_real=16'b0011111100100000; out_imag=16'b1111010101110010; end // in_theta = 1.947266 pi
 12'b111110010101: begin out_real=16'b0011111100100100; out_imag=16'b1111010110001011; end // in_theta = 1.947754 pi
 12'b111110010110: begin out_real=16'b0011111100101000; out_imag=16'b1111010110100100; end // in_theta = 1.948242 pi
 12'b111110010111: begin out_real=16'b0011111100101100; out_imag=16'b1111010110111100; end // in_theta = 1.948730 pi
 12'b111110011000: begin out_real=16'b0011111100110000; out_imag=16'b1111010111010101; end // in_theta = 1.949219 pi
 12'b111110011001: begin out_real=16'b0011111100110100; out_imag=16'b1111010111101110; end // in_theta = 1.949707 pi
 12'b111110011010: begin out_real=16'b0011111100111000; out_imag=16'b1111011000000111; end // in_theta = 1.950195 pi
 12'b111110011011: begin out_real=16'b0011111100111100; out_imag=16'b1111011000100000; end // in_theta = 1.950684 pi
 12'b111110011100: begin out_real=16'b0011111101000000; out_imag=16'b1111011000111001; end // in_theta = 1.951172 pi
 12'b111110011101: begin out_real=16'b0011111101000011; out_imag=16'b1111011001010001; end // in_theta = 1.951660 pi
 12'b111110011110: begin out_real=16'b0011111101000111; out_imag=16'b1111011001101010; end // in_theta = 1.952148 pi
 12'b111110011111: begin out_real=16'b0011111101001011; out_imag=16'b1111011010000011; end // in_theta = 1.952637 pi
 12'b111110100000: begin out_real=16'b0011111101001111; out_imag=16'b1111011010011100; end // in_theta = 1.953125 pi
 12'b111110100001: begin out_real=16'b0011111101010010; out_imag=16'b1111011010110101; end // in_theta = 1.953613 pi
 12'b111110100010: begin out_real=16'b0011111101010110; out_imag=16'b1111011011001110; end // in_theta = 1.954102 pi
 12'b111110100011: begin out_real=16'b0011111101011010; out_imag=16'b1111011011100111; end // in_theta = 1.954590 pi
 12'b111110100100: begin out_real=16'b0011111101011101; out_imag=16'b1111011011111111; end // in_theta = 1.955078 pi
 12'b111110100101: begin out_real=16'b0011111101100001; out_imag=16'b1111011100011000; end // in_theta = 1.955566 pi
 12'b111110100110: begin out_real=16'b0011111101100100; out_imag=16'b1111011100110001; end // in_theta = 1.956055 pi
 12'b111110100111: begin out_real=16'b0011111101101000; out_imag=16'b1111011101001010; end // in_theta = 1.956543 pi
 12'b111110101000: begin out_real=16'b0011111101101011; out_imag=16'b1111011101100011; end // in_theta = 1.957031 pi
 12'b111110101001: begin out_real=16'b0011111101101110; out_imag=16'b1111011101111100; end // in_theta = 1.957520 pi
 12'b111110101010: begin out_real=16'b0011111101110010; out_imag=16'b1111011110010101; end // in_theta = 1.958008 pi
 12'b111110101011: begin out_real=16'b0011111101110101; out_imag=16'b1111011110101110; end // in_theta = 1.958496 pi
 12'b111110101100: begin out_real=16'b0011111101111000; out_imag=16'b1111011111000111; end // in_theta = 1.958984 pi
 12'b111110101101: begin out_real=16'b0011111101111011; out_imag=16'b1111011111100000; end // in_theta = 1.959473 pi
 12'b111110101110: begin out_real=16'b0011111101111111; out_imag=16'b1111011111111001; end // in_theta = 1.959961 pi
 12'b111110101111: begin out_real=16'b0011111110000010; out_imag=16'b1111100000010001; end // in_theta = 1.960449 pi
 12'b111110110000: begin out_real=16'b0011111110000101; out_imag=16'b1111100000101010; end // in_theta = 1.960938 pi
 12'b111110110001: begin out_real=16'b0011111110001000; out_imag=16'b1111100001000011; end // in_theta = 1.961426 pi
 12'b111110110010: begin out_real=16'b0011111110001011; out_imag=16'b1111100001011100; end // in_theta = 1.961914 pi
 12'b111110110011: begin out_real=16'b0011111110001110; out_imag=16'b1111100001110101; end // in_theta = 1.962402 pi
 12'b111110110100: begin out_real=16'b0011111110010001; out_imag=16'b1111100010001110; end // in_theta = 1.962891 pi
 12'b111110110101: begin out_real=16'b0011111110010100; out_imag=16'b1111100010100111; end // in_theta = 1.963379 pi
 12'b111110110110: begin out_real=16'b0011111110010111; out_imag=16'b1111100011000000; end // in_theta = 1.963867 pi
 12'b111110110111: begin out_real=16'b0011111110011001; out_imag=16'b1111100011011001; end // in_theta = 1.964355 pi
 12'b111110111000: begin out_real=16'b0011111110011100; out_imag=16'b1111100011110010; end // in_theta = 1.964844 pi
 12'b111110111001: begin out_real=16'b0011111110011111; out_imag=16'b1111100100001011; end // in_theta = 1.965332 pi
 12'b111110111010: begin out_real=16'b0011111110100010; out_imag=16'b1111100100100100; end // in_theta = 1.965820 pi
 12'b111110111011: begin out_real=16'b0011111110100100; out_imag=16'b1111100100111101; end // in_theta = 1.966309 pi
 12'b111110111100: begin out_real=16'b0011111110100111; out_imag=16'b1111100101010110; end // in_theta = 1.966797 pi
 12'b111110111101: begin out_real=16'b0011111110101010; out_imag=16'b1111100101101111; end // in_theta = 1.967285 pi
 12'b111110111110: begin out_real=16'b0011111110101100; out_imag=16'b1111100110001000; end // in_theta = 1.967773 pi
 12'b111110111111: begin out_real=16'b0011111110101111; out_imag=16'b1111100110100001; end // in_theta = 1.968262 pi
 12'b111111000000: begin out_real=16'b0011111110110001; out_imag=16'b1111100110111010; end // in_theta = 1.968750 pi
 12'b111111000001: begin out_real=16'b0011111110110100; out_imag=16'b1111100111010011; end // in_theta = 1.969238 pi
 12'b111111000010: begin out_real=16'b0011111110110110; out_imag=16'b1111100111101100; end // in_theta = 1.969727 pi
 12'b111111000011: begin out_real=16'b0011111110111000; out_imag=16'b1111101000000101; end // in_theta = 1.970215 pi
 12'b111111000100: begin out_real=16'b0011111110111011; out_imag=16'b1111101000011110; end // in_theta = 1.970703 pi
 12'b111111000101: begin out_real=16'b0011111110111101; out_imag=16'b1111101000110111; end // in_theta = 1.971191 pi
 12'b111111000110: begin out_real=16'b0011111110111111; out_imag=16'b1111101001010000; end // in_theta = 1.971680 pi
 12'b111111000111: begin out_real=16'b0011111111000001; out_imag=16'b1111101001101001; end // in_theta = 1.972168 pi
 12'b111111001000: begin out_real=16'b0011111111000100; out_imag=16'b1111101010000010; end // in_theta = 1.972656 pi
 12'b111111001001: begin out_real=16'b0011111111000110; out_imag=16'b1111101010011011; end // in_theta = 1.973145 pi
 12'b111111001010: begin out_real=16'b0011111111001000; out_imag=16'b1111101010110100; end // in_theta = 1.973633 pi
 12'b111111001011: begin out_real=16'b0011111111001010; out_imag=16'b1111101011001101; end // in_theta = 1.974121 pi
 12'b111111001100: begin out_real=16'b0011111111001100; out_imag=16'b1111101011100110; end // in_theta = 1.974609 pi
 12'b111111001101: begin out_real=16'b0011111111001110; out_imag=16'b1111101100000000; end // in_theta = 1.975098 pi
 12'b111111001110: begin out_real=16'b0011111111010000; out_imag=16'b1111101100011001; end // in_theta = 1.975586 pi
 12'b111111001111: begin out_real=16'b0011111111010010; out_imag=16'b1111101100110010; end // in_theta = 1.976074 pi
 12'b111111010000: begin out_real=16'b0011111111010100; out_imag=16'b1111101101001011; end // in_theta = 1.976563 pi
 12'b111111010001: begin out_real=16'b0011111111010101; out_imag=16'b1111101101100100; end // in_theta = 1.977051 pi
 12'b111111010010: begin out_real=16'b0011111111010111; out_imag=16'b1111101101111101; end // in_theta = 1.977539 pi
 12'b111111010011: begin out_real=16'b0011111111011001; out_imag=16'b1111101110010110; end // in_theta = 1.978027 pi
 12'b111111010100: begin out_real=16'b0011111111011011; out_imag=16'b1111101110101111; end // in_theta = 1.978516 pi
 12'b111111010101: begin out_real=16'b0011111111011100; out_imag=16'b1111101111001000; end // in_theta = 1.979004 pi
 12'b111111010110: begin out_real=16'b0011111111011110; out_imag=16'b1111101111100001; end // in_theta = 1.979492 pi
 12'b111111010111: begin out_real=16'b0011111111100000; out_imag=16'b1111101111111010; end // in_theta = 1.979980 pi
 12'b111111011000: begin out_real=16'b0011111111100001; out_imag=16'b1111110000010011; end // in_theta = 1.980469 pi
 12'b111111011001: begin out_real=16'b0011111111100011; out_imag=16'b1111110000101100; end // in_theta = 1.980957 pi
 12'b111111011010: begin out_real=16'b0011111111100100; out_imag=16'b1111110001000101; end // in_theta = 1.981445 pi
 12'b111111011011: begin out_real=16'b0011111111100110; out_imag=16'b1111110001011111; end // in_theta = 1.981934 pi
 12'b111111011100: begin out_real=16'b0011111111100111; out_imag=16'b1111110001111000; end // in_theta = 1.982422 pi
 12'b111111011101: begin out_real=16'b0011111111101000; out_imag=16'b1111110010010001; end // in_theta = 1.982910 pi
 12'b111111011110: begin out_real=16'b0011111111101010; out_imag=16'b1111110010101010; end // in_theta = 1.983398 pi
 12'b111111011111: begin out_real=16'b0011111111101011; out_imag=16'b1111110011000011; end // in_theta = 1.983887 pi
 12'b111111100000: begin out_real=16'b0011111111101100; out_imag=16'b1111110011011100; end // in_theta = 1.984375 pi
 12'b111111100001: begin out_real=16'b0011111111101101; out_imag=16'b1111110011110101; end // in_theta = 1.984863 pi
 12'b111111100010: begin out_real=16'b0011111111101111; out_imag=16'b1111110100001110; end // in_theta = 1.985352 pi
 12'b111111100011: begin out_real=16'b0011111111110000; out_imag=16'b1111110100100111; end // in_theta = 1.985840 pi
 12'b111111100100: begin out_real=16'b0011111111110001; out_imag=16'b1111110101000000; end // in_theta = 1.986328 pi
 12'b111111100101: begin out_real=16'b0011111111110010; out_imag=16'b1111110101011010; end // in_theta = 1.986816 pi
 12'b111111100110: begin out_real=16'b0011111111110011; out_imag=16'b1111110101110011; end // in_theta = 1.987305 pi
 12'b111111100111: begin out_real=16'b0011111111110100; out_imag=16'b1111110110001100; end // in_theta = 1.987793 pi
 12'b111111101000: begin out_real=16'b0011111111110101; out_imag=16'b1111110110100101; end // in_theta = 1.988281 pi
 12'b111111101001: begin out_real=16'b0011111111110110; out_imag=16'b1111110110111110; end // in_theta = 1.988770 pi
 12'b111111101010: begin out_real=16'b0011111111110111; out_imag=16'b1111110111010111; end // in_theta = 1.989258 pi
 12'b111111101011: begin out_real=16'b0011111111110111; out_imag=16'b1111110111110000; end // in_theta = 1.989746 pi
 12'b111111101100: begin out_real=16'b0011111111111000; out_imag=16'b1111111000001001; end // in_theta = 1.990234 pi
 12'b111111101101: begin out_real=16'b0011111111111001; out_imag=16'b1111111000100011; end // in_theta = 1.990723 pi
 12'b111111101110: begin out_real=16'b0011111111111010; out_imag=16'b1111111000111100; end // in_theta = 1.991211 pi
 12'b111111101111: begin out_real=16'b0011111111111010; out_imag=16'b1111111001010101; end // in_theta = 1.991699 pi
 12'b111111110000: begin out_real=16'b0011111111111011; out_imag=16'b1111111001101110; end // in_theta = 1.992188 pi
 12'b111111110001: begin out_real=16'b0011111111111100; out_imag=16'b1111111010000111; end // in_theta = 1.992676 pi
 12'b111111110010: begin out_real=16'b0011111111111100; out_imag=16'b1111111010100000; end // in_theta = 1.993164 pi
 12'b111111110011: begin out_real=16'b0011111111111101; out_imag=16'b1111111010111001; end // in_theta = 1.993652 pi
 12'b111111110100: begin out_real=16'b0011111111111101; out_imag=16'b1111111011010010; end // in_theta = 1.994141 pi
 12'b111111110101: begin out_real=16'b0011111111111110; out_imag=16'b1111111011101100; end // in_theta = 1.994629 pi
 12'b111111110110: begin out_real=16'b0011111111111110; out_imag=16'b1111111100000101; end // in_theta = 1.995117 pi
 12'b111111110111: begin out_real=16'b0011111111111110; out_imag=16'b1111111100011110; end // in_theta = 1.995605 pi
 12'b111111111000: begin out_real=16'b0011111111111111; out_imag=16'b1111111100110111; end // in_theta = 1.996094 pi
 12'b111111111001: begin out_real=16'b0011111111111111; out_imag=16'b1111111101010000; end // in_theta = 1.996582 pi
 12'b111111111010: begin out_real=16'b0011111111111111; out_imag=16'b1111111101101001; end // in_theta = 1.997070 pi
 12'b111111111011: begin out_real=16'b0100000000000000; out_imag=16'b1111111110000010; end // in_theta = 1.997559 pi
 12'b111111111100: begin out_real=16'b0100000000000000; out_imag=16'b1111111110011011; end // in_theta = 1.998047 pi
 12'b111111111101: begin out_real=16'b0100000000000000; out_imag=16'b1111111110110101; end // in_theta = 1.998535 pi
 12'b111111111110: begin out_real=16'b0100000000000000; out_imag=16'b1111111111001110; end // in_theta = 1.999023 pi
 12'b111111111111: begin out_real=16'b0100000000000000; out_imag=16'b1111111111100111; end // in_theta = 1.999512 pi
 endcase
end
endmodule
