module adder_5bit_11_tb();
reg [4:0] in0;
reg [4:0] in1;
reg [4:0] in2;
reg [4:0] in3;
reg [4:0] in4;
reg [4:0] in5;
reg [4:0] in6;
reg [4:0] in7;
reg [4:0] in8;
reg [4:0] in9;
reg [4:0] in10;
wire [4:0] out;

adder_5bit_11 testbench_instatiation(in0[4:0],in1[4:0],in2[4:0],in3[4:0],in4[4:0],in5[4:0],in6[4:0],in7[4:0],in8[4:0],in9[4:0],in10[4:0],out[4:0]);

initial begin
$monitor($time,"out=%b",out[4:0]);
# 10;
in0[4:0]=5'b10101;
in1[4:0]=5'b10101;
in2[4:0]=5'b10101;
in3[4:0]=5'b10101;
in4[4:0]=5'b10101;
in5[4:0]=5'b10101;
in6[4:0]=5'b10101;
in7[4:0]=5'b10101;
in8[4:0]=5'b10101;
in9[4:0]=5'b10101;
in10[4:0]=5'b10101;
# 50;
in0[4:0]=5'b11101;
in1[4:0]=5'b11101;
in2[4:0]=5'b11101;
in3[4:0]=5'b11101;
in4[4:0]=5'b11101;
in5[4:0]=5'b11101;
in6[4:0]=5'b11101;
in7[4:0]=5'b11101;
in8[4:0]=5'b11101;
in9[4:0]=5'b11101;
in10[4:0]=5'b11101;
# 50;
end
endmodule
