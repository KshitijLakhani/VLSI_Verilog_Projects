module FFT (
input clk,
input reg [11:0] wn_exp,            //theta
input reg [15:0] a_r,                  
input reg [15:0] a_i,
input reg [15:0] b_r,                  
input reg [15:0] b_i,
output reg [15:0] x_r,            
output reg [15:0] x_i,
output reg [15:0] y_r,
output reg [15:0] y_i);

// Declarations for sequential part
reg [15:0] wn_exp_out;
reg [15:0] a_r_out;                  
reg [15:0] a_i_out;
reg [15:0] b_r_out;                 
reg [15:0] b_i_out;


// Declarations for Wn 
wire [15:0] realout;
wire [15:0] imagout;


//Extra Declarations for Xgen and Ygen
/*reg [15:0] x_real_reg;
reg [15:0] x_imag_reg;
reg [15:0] y_real_reg;
reg [15:0] y_imag_reg;*/

// Declarations for Xgen and Ygen
wire [15:0] x_real;
wire [15:0] x_imag;
wire [15:0] y_real;
wire [15:0] y_imag;


//Sequential part 
always@(posedge clk)begin
// Making all the inputs change on positive clock edge only
wn_exp_out <= #1 wn_exp;
a_r_out <= #1 a_r;
a_i_out <= #1 a_i;
b_r_out <= #1 b_r;
b_i_out <= #1 b_i;

// Actual outputs being assigned on positive clock edge only

x_r <= #1 x_real;
x_i <= #1 x_imag;
y_r <= #1 y_real;
y_i <= #1 y_imag;

end


Wngenerator Wngen(clk,wn_exp,realout,imagout);
Xgenerator Xgen(a_r_out,a_i_out,b_r_out,b_i_out,x_real,x_imag);
Ygenerator Ygen(a_r_out,a_i_out,b_r_out,b_i_out,realout,imagout,y_real,y_imag);

endmodule



// X generator
module Xgenerator (
input [15:0] a_re,
input [15:0] a_im,
input [15:0] b_re,
input [15:0] b_im,
output reg [15:0] x_real,
output reg [15:0] x_imag);

always @ (a_re or a_im or b_im or b_re) begin
x_real=a_re + b_re;
x_imag=a_im + b_im;
end

endmodule

// Y generator
module Ygenerator (
input [15:0] a_re,
input [15:0] a_im,
input [15:0] b_re,
input [15:0] b_im,
input [15:0] w_r,
input [15:0] w_i,
output reg [15:0] y_real,
output reg [15:0] y_imag);

reg [16:0] temp_r_r;
reg [16:0] temp_i_i;
reg [32:0] temp_r;
reg [32:0] temp_i;

always @ (a_re or a_im or b_im or b_re or w_r or w_i) begin

//(A-B)- 17 bits
temp_r_r=a_re - b_re;
temp_i_i=a_im - b_im;
//(A-B)*Wn - 33 bits
temp_r=(temp_r_r)*(w_r) - (temp_i_i)*(w_i);
temp_i=(temp_i_i)*(w_r) - (temp_r_r)*(w_i);
//(A-B)*Wn - 16 bits
y_real=temp_r[32:17];
y_imag=temp_i[32:17];
end
endmodule
// Wn gen
module Wngenerator(
input clk,
input [11:0] in_theta,
output reg [15:0]realout,
output reg [15:0]imagout);


//wire [11:0]in_theta;
//wire clk;
//reg [15:0]realout;
//reg [15:0]imagout;

reg [11:0]theta;
reg [11:0]thegen1;
reg [11:0]thegen;
reg [15:0]real3;
reg [15:0]imag3;
reg [15:0]real2;
reg [15:0]imag2;
reg [15:0]real1;
reg [15:0]imag1;
reg [15:0]tmp;

always@(posedge clk)begin
theta<= #1 in_theta;
realout<= #1 real3;
imagout<= #1 imag3;
end

always @(*) begin
if (theta<=12'b010000000000)begin
    thegen = theta;
    real3 =real1;
    imag3=imag1; end
else if (theta<=12'b100000000000 && theta>12'b010000000000)begin
    thegen = 12'b100000000000-theta;
    real3 =~real1+1'b1;
    imag3=imag1; end
else if (theta<=12'b110000000000 && theta>12'b100000000000)begin
    thegen = theta-12'b100000000000;
    real3 = ~real1+1'b1;
    imag3=~imag1+1'b1; end
else if (theta<=12'b111111111111 && theta>12'b110000000000)begin
    thegen = 12'b111111111111-theta+1'b1;
    real3 = real1;
    imag3=~imag1+1'b1; end
end
always @(*)begin
if (thegen>12'b001000000000)begin
    thegen1=12'b010000000000-thegen;
    tmp=imag1;    
    imag1=real1;    
    real1=tmp;
end
else if(thegen<=12'b001000000000)begin
    thegen1=thegen;
end
end

always @(thegen1) begin
  case (thegen1)
    12'b000000000000: begin  real1=16'b0100000000000000; imag1=16'b0000000000000000;  end  // angle = 0.000000 pi
    12'b000000000001: begin  real1=16'b0100000000000000; imag1=16'b0000000000011001;  end  // angle = 0.000488 pi
    12'b000000000010: begin  real1=16'b0100000000000000; imag1=16'b0000000000110010;  end  // angle = 0.000977 pi
    12'b000000000011: begin  real1=16'b0100000000000000; imag1=16'b0000000001001011;  end  // angle = 0.001465 pi
    12'b000000000100: begin  real1=16'b0100000000000000; imag1=16'b0000000001100101;  end  // angle = 0.001953 pi
    12'b000000000101: begin  real1=16'b0100000000000000; imag1=16'b0000000001111110;  end  // angle = 0.002441 pi
    12'b000000000110: begin  real1=16'b0011111111111111; imag1=16'b0000000010010111;  end  // angle = 0.002930 pi
    12'b000000000111: begin  real1=16'b0011111111111111; imag1=16'b0000000010110000;  end  // angle = 0.003418 pi
    12'b000000001000: begin  real1=16'b0011111111111111; imag1=16'b0000000011001001;  end  // angle = 0.003906 pi
    12'b000000001001: begin  real1=16'b0011111111111110; imag1=16'b0000000011100010;  end  // angle = 0.004395 pi
    12'b000000001010: begin  real1=16'b0011111111111110; imag1=16'b0000000011111011;  end  // angle = 0.004883 pi
    12'b000000001011: begin  real1=16'b0011111111111110; imag1=16'b0000000100010100;  end  // angle = 0.005371 pi
    12'b000000001100: begin  real1=16'b0011111111111101; imag1=16'b0000000100101110;  end  // angle = 0.005859 pi
    12'b000000001101: begin  real1=16'b0011111111111101; imag1=16'b0000000101000111;  end  // angle = 0.006348 pi
    12'b000000001110: begin  real1=16'b0011111111111100; imag1=16'b0000000101100000;  end  // angle = 0.006836 pi
    12'b000000001111: begin  real1=16'b0011111111111100; imag1=16'b0000000101111001;  end  // angle = 0.007324 pi
    12'b000000010000: begin  real1=16'b0011111111111011; imag1=16'b0000000110010010;  end  // angle = 0.007812 pi
    12'b000000010001: begin  real1=16'b0011111111111010; imag1=16'b0000000110101011;  end  // angle = 0.008301 pi
    12'b000000010010: begin  real1=16'b0011111111111010; imag1=16'b0000000111000100;  end  // angle = 0.008789 pi
    12'b000000010011: begin  real1=16'b0011111111111001; imag1=16'b0000000111011101;  end  // angle = 0.009277 pi
    12'b000000010100: begin  real1=16'b0011111111111000; imag1=16'b0000000111110111;  end  // angle = 0.009766 pi
    12'b000000010101: begin  real1=16'b0011111111110111; imag1=16'b0000001000010000;  end  // angle = 0.010254 pi
    12'b000000010110: begin  real1=16'b0011111111110111; imag1=16'b0000001000101001;  end  // angle = 0.010742 pi
    12'b000000010111: begin  real1=16'b0011111111110110; imag1=16'b0000001001000010;  end  // angle = 0.011230 pi
    12'b000000011000: begin  real1=16'b0011111111110101; imag1=16'b0000001001011011;  end  // angle = 0.011719 pi
    12'b000000011001: begin  real1=16'b0011111111110100; imag1=16'b0000001001110100;  end  // angle = 0.012207 pi
    12'b000000011010: begin  real1=16'b0011111111110011; imag1=16'b0000001010001101;  end  // angle = 0.012695 pi
    12'b000000011011: begin  real1=16'b0011111111110010; imag1=16'b0000001010100110;  end  // angle = 0.013184 pi
    12'b000000011100: begin  real1=16'b0011111111110001; imag1=16'b0000001011000000;  end  // angle = 0.013672 pi
    12'b000000011101: begin  real1=16'b0011111111110000; imag1=16'b0000001011011001;  end  // angle = 0.014160 pi
    12'b000000011110: begin  real1=16'b0011111111101111; imag1=16'b0000001011110010;  end  // angle = 0.014648 pi
    12'b000000011111: begin  real1=16'b0011111111101101; imag1=16'b0000001100001011;  end  // angle = 0.015137 pi
    12'b000000100000: begin  real1=16'b0011111111101100; imag1=16'b0000001100100100;  end  // angle = 0.015625 pi
    12'b000000100001: begin  real1=16'b0011111111101011; imag1=16'b0000001100111101;  end  // angle = 0.016113 pi
    12'b000000100010: begin  real1=16'b0011111111101010; imag1=16'b0000001101010110;  end  // angle = 0.016602 pi
    12'b000000100011: begin  real1=16'b0011111111101000; imag1=16'b0000001101101111;  end  // angle = 0.017090 pi
    12'b000000100100: begin  real1=16'b0011111111100111; imag1=16'b0000001110001000;  end  // angle = 0.017578 pi
    12'b000000100101: begin  real1=16'b0011111111100110; imag1=16'b0000001110100001;  end  // angle = 0.018066 pi
    12'b000000100110: begin  real1=16'b0011111111100100; imag1=16'b0000001110111011;  end  // angle = 0.018555 pi
    12'b000000100111: begin  real1=16'b0011111111100011; imag1=16'b0000001111010100;  end  // angle = 0.019043 pi
    12'b000000101000: begin  real1=16'b0011111111100001; imag1=16'b0000001111101101;  end  // angle = 0.019531 pi
    12'b000000101001: begin  real1=16'b0011111111100000; imag1=16'b0000010000000110;  end  // angle = 0.020020 pi
    12'b000000101010: begin  real1=16'b0011111111011110; imag1=16'b0000010000011111;  end  // angle = 0.020508 pi
    12'b000000101011: begin  real1=16'b0011111111011100; imag1=16'b0000010000111000;  end  // angle = 0.020996 pi
    12'b000000101100: begin  real1=16'b0011111111011011; imag1=16'b0000010001010001;  end  // angle = 0.021484 pi
    12'b000000101101: begin  real1=16'b0011111111011001; imag1=16'b0000010001101010;  end  // angle = 0.021973 pi
    12'b000000101110: begin  real1=16'b0011111111010111; imag1=16'b0000010010000011;  end  // angle = 0.022461 pi
    12'b000000101111: begin  real1=16'b0011111111010101; imag1=16'b0000010010011100;  end  // angle = 0.022949 pi
    12'b000000110000: begin  real1=16'b0011111111010100; imag1=16'b0000010010110101;  end  // angle = 0.023438 pi
    12'b000000110001: begin  real1=16'b0011111111010010; imag1=16'b0000010011001110;  end  // angle = 0.023926 pi
    12'b000000110010: begin  real1=16'b0011111111010000; imag1=16'b0000010011100111;  end  // angle = 0.024414 pi
    12'b000000110011: begin  real1=16'b0011111111001110; imag1=16'b0000010100000000;  end  // angle = 0.024902 pi
    12'b000000110100: begin  real1=16'b0011111111001100; imag1=16'b0000010100011010;  end  // angle = 0.025391 pi
    12'b000000110101: begin  real1=16'b0011111111001010; imag1=16'b0000010100110011;  end  // angle = 0.025879 pi
    12'b000000110110: begin  real1=16'b0011111111001000; imag1=16'b0000010101001100;  end  // angle = 0.026367 pi
    12'b000000110111: begin  real1=16'b0011111111000110; imag1=16'b0000010101100101;  end  // angle = 0.026855 pi
    12'b000000111000: begin  real1=16'b0011111111000100; imag1=16'b0000010101111110;  end  // angle = 0.027344 pi
    12'b000000111001: begin  real1=16'b0011111111000001; imag1=16'b0000010110010111;  end  // angle = 0.027832 pi
    12'b000000111010: begin  real1=16'b0011111110111111; imag1=16'b0000010110110000;  end  // angle = 0.028320 pi
    12'b000000111011: begin  real1=16'b0011111110111101; imag1=16'b0000010111001001;  end  // angle = 0.028809 pi
    12'b000000111100: begin  real1=16'b0011111110111011; imag1=16'b0000010111100010;  end  // angle = 0.029297 pi
    12'b000000111101: begin  real1=16'b0011111110111000; imag1=16'b0000010111111011;  end  // angle = 0.029785 pi
    12'b000000111110: begin  real1=16'b0011111110110110; imag1=16'b0000011000010100;  end  // angle = 0.030273 pi
    12'b000000111111: begin  real1=16'b0011111110110100; imag1=16'b0000011000101101;  end  // angle = 0.030762 pi
    12'b000001000000: begin  real1=16'b0011111110110001; imag1=16'b0000011001000110;  end  // angle = 0.031250 pi
    12'b000001000001: begin  real1=16'b0011111110101111; imag1=16'b0000011001011111;  end  // angle = 0.031738 pi
    12'b000001000010: begin  real1=16'b0011111110101100; imag1=16'b0000011001111000;  end  // angle = 0.032227 pi
    12'b000001000011: begin  real1=16'b0011111110101010; imag1=16'b0000011010010001;  end  // angle = 0.032715 pi
    12'b000001000100: begin  real1=16'b0011111110100111; imag1=16'b0000011010101010;  end  // angle = 0.033203 pi
    12'b000001000101: begin  real1=16'b0011111110100100; imag1=16'b0000011011000011;  end  // angle = 0.033691 pi
    12'b000001000110: begin  real1=16'b0011111110100010; imag1=16'b0000011011011100;  end  // angle = 0.034180 pi
    12'b000001000111: begin  real1=16'b0011111110011111; imag1=16'b0000011011110101;  end  // angle = 0.034668 pi
    12'b000001001000: begin  real1=16'b0011111110011100; imag1=16'b0000011100001110;  end  // angle = 0.035156 pi
    12'b000001001001: begin  real1=16'b0011111110011001; imag1=16'b0000011100100111;  end  // angle = 0.035645 pi
    12'b000001001010: begin  real1=16'b0011111110010111; imag1=16'b0000011101000000;  end  // angle = 0.036133 pi
    12'b000001001011: begin  real1=16'b0011111110010100; imag1=16'b0000011101011001;  end  // angle = 0.036621 pi
    12'b000001001100: begin  real1=16'b0011111110010001; imag1=16'b0000011101110010;  end  // angle = 0.037109 pi
    12'b000001001101: begin  real1=16'b0011111110001110; imag1=16'b0000011110001011;  end  // angle = 0.037598 pi
    12'b000001001110: begin  real1=16'b0011111110001011; imag1=16'b0000011110100100;  end  // angle = 0.038086 pi
    12'b000001001111: begin  real1=16'b0011111110001000; imag1=16'b0000011110111101;  end  // angle = 0.038574 pi
    12'b000001010000: begin  real1=16'b0011111110000101; imag1=16'b0000011111010110;  end  // angle = 0.039062 pi
    12'b000001010001: begin  real1=16'b0011111110000010; imag1=16'b0000011111101111;  end  // angle = 0.039551 pi
    12'b000001010010: begin  real1=16'b0011111101111111; imag1=16'b0000100000000111;  end  // angle = 0.040039 pi
    12'b000001010011: begin  real1=16'b0011111101111011; imag1=16'b0000100000100000;  end  // angle = 0.040527 pi
    12'b000001010100: begin  real1=16'b0011111101111000; imag1=16'b0000100000111001;  end  // angle = 0.041016 pi
    12'b000001010101: begin  real1=16'b0011111101110101; imag1=16'b0000100001010010;  end  // angle = 0.041504 pi
    12'b000001010110: begin  real1=16'b0011111101110010; imag1=16'b0000100001101011;  end  // angle = 0.041992 pi
    12'b000001010111: begin  real1=16'b0011111101101110; imag1=16'b0000100010000100;  end  // angle = 0.042480 pi
    12'b000001011000: begin  real1=16'b0011111101101011; imag1=16'b0000100010011101;  end  // angle = 0.042969 pi
    12'b000001011001: begin  real1=16'b0011111101101000; imag1=16'b0000100010110110;  end  // angle = 0.043457 pi
    12'b000001011010: begin  real1=16'b0011111101100100; imag1=16'b0000100011001111;  end  // angle = 0.043945 pi
    12'b000001011011: begin  real1=16'b0011111101100001; imag1=16'b0000100011101000;  end  // angle = 0.044434 pi
    12'b000001011100: begin  real1=16'b0011111101011101; imag1=16'b0000100100000001;  end  // angle = 0.044922 pi
    12'b000001011101: begin  real1=16'b0011111101011010; imag1=16'b0000100100011001;  end  // angle = 0.045410 pi
    12'b000001011110: begin  real1=16'b0011111101010110; imag1=16'b0000100100110010;  end  // angle = 0.045898 pi
    12'b000001011111: begin  real1=16'b0011111101010010; imag1=16'b0000100101001011;  end  // angle = 0.046387 pi
    12'b000001100000: begin  real1=16'b0011111101001111; imag1=16'b0000100101100100;  end  // angle = 0.046875 pi
    12'b000001100001: begin  real1=16'b0011111101001011; imag1=16'b0000100101111101;  end  // angle = 0.047363 pi
    12'b000001100010: begin  real1=16'b0011111101000111; imag1=16'b0000100110010110;  end  // angle = 0.047852 pi
    12'b000001100011: begin  real1=16'b0011111101000011; imag1=16'b0000100110101111;  end  // angle = 0.048340 pi
    12'b000001100100: begin  real1=16'b0011111101000000; imag1=16'b0000100111000111;  end  // angle = 0.048828 pi
    12'b000001100101: begin  real1=16'b0011111100111100; imag1=16'b0000100111100000;  end  // angle = 0.049316 pi
    12'b000001100110: begin  real1=16'b0011111100111000; imag1=16'b0000100111111001;  end  // angle = 0.049805 pi
    12'b000001100111: begin  real1=16'b0011111100110100; imag1=16'b0000101000010010;  end  // angle = 0.050293 pi
    12'b000001101000: begin  real1=16'b0011111100110000; imag1=16'b0000101000101011;  end  // angle = 0.050781 pi
    12'b000001101001: begin  real1=16'b0011111100101100; imag1=16'b0000101001000100;  end  // angle = 0.051270 pi
    12'b000001101010: begin  real1=16'b0011111100101000; imag1=16'b0000101001011100;  end  // angle = 0.051758 pi
    12'b000001101011: begin  real1=16'b0011111100100100; imag1=16'b0000101001110101;  end  // angle = 0.052246 pi
    12'b000001101100: begin  real1=16'b0011111100100000; imag1=16'b0000101010001110;  end  // angle = 0.052734 pi
    12'b000001101101: begin  real1=16'b0011111100011100; imag1=16'b0000101010100111;  end  // angle = 0.053223 pi
    12'b000001101110: begin  real1=16'b0011111100010111; imag1=16'b0000101011000000;  end  // angle = 0.053711 pi
    12'b000001101111: begin  real1=16'b0011111100010011; imag1=16'b0000101011011000;  end  // angle = 0.054199 pi
    12'b000001110000: begin  real1=16'b0011111100001111; imag1=16'b0000101011110001;  end  // angle = 0.054688 pi
    12'b000001110001: begin  real1=16'b0011111100001010; imag1=16'b0000101100001010;  end  // angle = 0.055176 pi
    12'b000001110010: begin  real1=16'b0011111100000110; imag1=16'b0000101100100011;  end  // angle = 0.055664 pi
    12'b000001110011: begin  real1=16'b0011111100000010; imag1=16'b0000101100111011;  end  // angle = 0.056152 pi
    12'b000001110100: begin  real1=16'b0011111011111101; imag1=16'b0000101101010100;  end  // angle = 0.056641 pi
    12'b000001110101: begin  real1=16'b0011111011111001; imag1=16'b0000101101101101;  end  // angle = 0.057129 pi
    12'b000001110110: begin  real1=16'b0011111011110100; imag1=16'b0000101110000101;  end  // angle = 0.057617 pi
    12'b000001110111: begin  real1=16'b0011111011110000; imag1=16'b0000101110011110;  end  // angle = 0.058105 pi
    12'b000001111000: begin  real1=16'b0011111011101011; imag1=16'b0000101110110111;  end  // angle = 0.058594 pi
    12'b000001111001: begin  real1=16'b0011111011100111; imag1=16'b0000101111010000;  end  // angle = 0.059082 pi
    12'b000001111010: begin  real1=16'b0011111011100010; imag1=16'b0000101111101000;  end  // angle = 0.059570 pi
    12'b000001111011: begin  real1=16'b0011111011011101; imag1=16'b0000110000000001;  end  // angle = 0.060059 pi
    12'b000001111100: begin  real1=16'b0011111011011000; imag1=16'b0000110000011010;  end  // angle = 0.060547 pi
    12'b000001111101: begin  real1=16'b0011111011010100; imag1=16'b0000110000110010;  end  // angle = 0.061035 pi
    12'b000001111110: begin  real1=16'b0011111011001111; imag1=16'b0000110001001011;  end  // angle = 0.061523 pi
    12'b000001111111: begin  real1=16'b0011111011001010; imag1=16'b0000110001100100;  end  // angle = 0.062012 pi
    12'b000010000000: begin  real1=16'b0011111011000101; imag1=16'b0000110001111100;  end  // angle = 0.062500 pi
    12'b000010000001: begin  real1=16'b0011111011000000; imag1=16'b0000110010010101;  end  // angle = 0.062988 pi
    12'b000010000010: begin  real1=16'b0011111010111011; imag1=16'b0000110010101110;  end  // angle = 0.063477 pi
    12'b000010000011: begin  real1=16'b0011111010110110; imag1=16'b0000110011000110;  end  // angle = 0.063965 pi
    12'b000010000100: begin  real1=16'b0011111010110001; imag1=16'b0000110011011111;  end  // angle = 0.064453 pi
    12'b000010000101: begin  real1=16'b0011111010101100; imag1=16'b0000110011111000;  end  // angle = 0.064941 pi
    12'b000010000110: begin  real1=16'b0011111010100111; imag1=16'b0000110100010000;  end  // angle = 0.065430 pi
    12'b000010000111: begin  real1=16'b0011111010100010; imag1=16'b0000110100101001;  end  // angle = 0.065918 pi
    12'b000010001000: begin  real1=16'b0011111010011101; imag1=16'b0000110101000001;  end  // angle = 0.066406 pi
    12'b000010001001: begin  real1=16'b0011111010011000; imag1=16'b0000110101011010;  end  // angle = 0.066895 pi
    12'b000010001010: begin  real1=16'b0011111010010010; imag1=16'b0000110101110010;  end  // angle = 0.067383 pi
    12'b000010001011: begin  real1=16'b0011111010001101; imag1=16'b0000110110001011;  end  // angle = 0.067871 pi
    12'b000010001100: begin  real1=16'b0011111010001000; imag1=16'b0000110110100100;  end  // angle = 0.068359 pi
    12'b000010001101: begin  real1=16'b0011111010000010; imag1=16'b0000110110111100;  end  // angle = 0.068848 pi
    12'b000010001110: begin  real1=16'b0011111001111101; imag1=16'b0000110111010101;  end  // angle = 0.069336 pi
    12'b000010001111: begin  real1=16'b0011111001110111; imag1=16'b0000110111101101;  end  // angle = 0.069824 pi
    12'b000010010000: begin  real1=16'b0011111001110010; imag1=16'b0000111000000110;  end  // angle = 0.070312 pi
    12'b000010010001: begin  real1=16'b0011111001101100; imag1=16'b0000111000011110;  end  // angle = 0.070801 pi
    12'b000010010010: begin  real1=16'b0011111001100111; imag1=16'b0000111000110111;  end  // angle = 0.071289 pi
    12'b000010010011: begin  real1=16'b0011111001100001; imag1=16'b0000111001001111;  end  // angle = 0.071777 pi
    12'b000010010100: begin  real1=16'b0011111001011100; imag1=16'b0000111001101000;  end  // angle = 0.072266 pi
    12'b000010010101: begin  real1=16'b0011111001010110; imag1=16'b0000111010000000;  end  // angle = 0.072754 pi
    12'b000010010110: begin  real1=16'b0011111001010000; imag1=16'b0000111010011001;  end  // angle = 0.073242 pi
    12'b000010010111: begin  real1=16'b0011111001001010; imag1=16'b0000111010110001;  end  // angle = 0.073730 pi
    12'b000010011000: begin  real1=16'b0011111001000101; imag1=16'b0000111011001010;  end  // angle = 0.074219 pi
    12'b000010011001: begin  real1=16'b0011111000111111; imag1=16'b0000111011100010;  end  // angle = 0.074707 pi
    12'b000010011010: begin  real1=16'b0011111000111001; imag1=16'b0000111011111011;  end  // angle = 0.075195 pi
    12'b000010011011: begin  real1=16'b0011111000110011; imag1=16'b0000111100010011;  end  // angle = 0.075684 pi
    12'b000010011100: begin  real1=16'b0011111000101101; imag1=16'b0000111100101011;  end  // angle = 0.076172 pi
    12'b000010011101: begin  real1=16'b0011111000100111; imag1=16'b0000111101000100;  end  // angle = 0.076660 pi
    12'b000010011110: begin  real1=16'b0011111000100001; imag1=16'b0000111101011100;  end  // angle = 0.077148 pi
    12'b000010011111: begin  real1=16'b0011111000011011; imag1=16'b0000111101110101;  end  // angle = 0.077637 pi
    12'b000010100000: begin  real1=16'b0011111000010101; imag1=16'b0000111110001101;  end  // angle = 0.078125 pi
    12'b000010100001: begin  real1=16'b0011111000001111; imag1=16'b0000111110100101;  end  // angle = 0.078613 pi
    12'b000010100010: begin  real1=16'b0011111000001001; imag1=16'b0000111110111110;  end  // angle = 0.079102 pi
    12'b000010100011: begin  real1=16'b0011111000000011; imag1=16'b0000111111010110;  end  // angle = 0.079590 pi
    12'b000010100100: begin  real1=16'b0011110111111100; imag1=16'b0000111111101110;  end  // angle = 0.080078 pi
    12'b000010100101: begin  real1=16'b0011110111110110; imag1=16'b0001000000000111;  end  // angle = 0.080566 pi
    12'b000010100110: begin  real1=16'b0011110111110000; imag1=16'b0001000000011111;  end  // angle = 0.081055 pi
    12'b000010100111: begin  real1=16'b0011110111101001; imag1=16'b0001000000110111;  end  // angle = 0.081543 pi
    12'b000010101000: begin  real1=16'b0011110111100011; imag1=16'b0001000001010000;  end  // angle = 0.082031 pi
    12'b000010101001: begin  real1=16'b0011110111011101; imag1=16'b0001000001101000;  end  // angle = 0.082520 pi
    12'b000010101010: begin  real1=16'b0011110111010110; imag1=16'b0001000010000000;  end  // angle = 0.083008 pi
    12'b000010101011: begin  real1=16'b0011110111010000; imag1=16'b0001000010011001;  end  // angle = 0.083496 pi
    12'b000010101100: begin  real1=16'b0011110111001001; imag1=16'b0001000010110001;  end  // angle = 0.083984 pi
    12'b000010101101: begin  real1=16'b0011110111000010; imag1=16'b0001000011001001;  end  // angle = 0.084473 pi
    12'b000010101110: begin  real1=16'b0011110110111100; imag1=16'b0001000011100001;  end  // angle = 0.084961 pi
    12'b000010101111: begin  real1=16'b0011110110110101; imag1=16'b0001000011111010;  end  // angle = 0.085449 pi
    12'b000010110000: begin  real1=16'b0011110110101111; imag1=16'b0001000100010010;  end  // angle = 0.085937 pi
    12'b000010110001: begin  real1=16'b0011110110101000; imag1=16'b0001000100101010;  end  // angle = 0.086426 pi
    12'b000010110010: begin  real1=16'b0011110110100001; imag1=16'b0001000101000010;  end  // angle = 0.086914 pi
    12'b000010110011: begin  real1=16'b0011110110011010; imag1=16'b0001000101011010;  end  // angle = 0.087402 pi
    12'b000010110100: begin  real1=16'b0011110110010011; imag1=16'b0001000101110011;  end  // angle = 0.087891 pi
    12'b000010110101: begin  real1=16'b0011110110001101; imag1=16'b0001000110001011;  end  // angle = 0.088379 pi
    12'b000010110110: begin  real1=16'b0011110110000110; imag1=16'b0001000110100011;  end  // angle = 0.088867 pi
    12'b000010110111: begin  real1=16'b0011110101111111; imag1=16'b0001000110111011;  end  // angle = 0.089355 pi
    12'b000010111000: begin  real1=16'b0011110101111000; imag1=16'b0001000111010011;  end  // angle = 0.089844 pi
    12'b000010111001: begin  real1=16'b0011110101110001; imag1=16'b0001000111101011;  end  // angle = 0.090332 pi
    12'b000010111010: begin  real1=16'b0011110101101010; imag1=16'b0001001000000100;  end  // angle = 0.090820 pi
    12'b000010111011: begin  real1=16'b0011110101100011; imag1=16'b0001001000011100;  end  // angle = 0.091309 pi
    12'b000010111100: begin  real1=16'b0011110101011011; imag1=16'b0001001000110100;  end  // angle = 0.091797 pi
    12'b000010111101: begin  real1=16'b0011110101010100; imag1=16'b0001001001001100;  end  // angle = 0.092285 pi
    12'b000010111110: begin  real1=16'b0011110101001101; imag1=16'b0001001001100100;  end  // angle = 0.092773 pi
    12'b000010111111: begin  real1=16'b0011110101000110; imag1=16'b0001001001111100;  end  // angle = 0.093262 pi
    12'b000011000000: begin  real1=16'b0011110100111111; imag1=16'b0001001010010100;  end  // angle = 0.093750 pi
    12'b000011000001: begin  real1=16'b0011110100110111; imag1=16'b0001001010101100;  end  // angle = 0.094238 pi
    12'b000011000010: begin  real1=16'b0011110100110000; imag1=16'b0001001011000100;  end  // angle = 0.094727 pi
    12'b000011000011: begin  real1=16'b0011110100101000; imag1=16'b0001001011011100;  end  // angle = 0.095215 pi
    12'b000011000100: begin  real1=16'b0011110100100001; imag1=16'b0001001011110100;  end  // angle = 0.095703 pi
    12'b000011000101: begin  real1=16'b0011110100011010; imag1=16'b0001001100001100;  end  // angle = 0.096191 pi
    12'b000011000110: begin  real1=16'b0011110100010010; imag1=16'b0001001100100100;  end  // angle = 0.096680 pi
    12'b000011000111: begin  real1=16'b0011110100001011; imag1=16'b0001001100111100;  end  // angle = 0.097168 pi
    12'b000011001000: begin  real1=16'b0011110100000011; imag1=16'b0001001101010100;  end  // angle = 0.097656 pi
    12'b000011001001: begin  real1=16'b0011110011111011; imag1=16'b0001001101101100;  end  // angle = 0.098145 pi
    12'b000011001010: begin  real1=16'b0011110011110100; imag1=16'b0001001110000100;  end  // angle = 0.098633 pi
    12'b000011001011: begin  real1=16'b0011110011101100; imag1=16'b0001001110011100;  end  // angle = 0.099121 pi
    12'b000011001100: begin  real1=16'b0011110011100100; imag1=16'b0001001110110100;  end  // angle = 0.099609 pi
    12'b000011001101: begin  real1=16'b0011110011011101; imag1=16'b0001001111001100;  end  // angle = 0.100098 pi
    12'b000011001110: begin  real1=16'b0011110011010101; imag1=16'b0001001111100100;  end  // angle = 0.100586 pi
    12'b000011001111: begin  real1=16'b0011110011001101; imag1=16'b0001001111111011;  end  // angle = 0.101074 pi
    12'b000011010000: begin  real1=16'b0011110011000101; imag1=16'b0001010000010011;  end  // angle = 0.101563 pi
    12'b000011010001: begin  real1=16'b0011110010111101; imag1=16'b0001010000101011;  end  // angle = 0.102051 pi
    12'b000011010010: begin  real1=16'b0011110010110101; imag1=16'b0001010001000011;  end  // angle = 0.102539 pi
    12'b000011010011: begin  real1=16'b0011110010101101; imag1=16'b0001010001011011;  end  // angle = 0.103027 pi
    12'b000011010100: begin  real1=16'b0011110010100101; imag1=16'b0001010001110011;  end  // angle = 0.103516 pi
    12'b000011010101: begin  real1=16'b0011110010011101; imag1=16'b0001010010001011;  end  // angle = 0.104004 pi
    12'b000011010110: begin  real1=16'b0011110010010101; imag1=16'b0001010010100010;  end  // angle = 0.104492 pi
    12'b000011010111: begin  real1=16'b0011110010001101; imag1=16'b0001010010111010;  end  // angle = 0.104980 pi
    12'b000011011000: begin  real1=16'b0011110010000101; imag1=16'b0001010011010010;  end  // angle = 0.105469 pi
    12'b000011011001: begin  real1=16'b0011110001111101; imag1=16'b0001010011101010;  end  // angle = 0.105957 pi
    12'b000011011010: begin  real1=16'b0011110001110100; imag1=16'b0001010100000001;  end  // angle = 0.106445 pi
    12'b000011011011: begin  real1=16'b0011110001101100; imag1=16'b0001010100011001;  end  // angle = 0.106934 pi
    12'b000011011100: begin  real1=16'b0011110001100100; imag1=16'b0001010100110001;  end  // angle = 0.107422 pi
    12'b000011011101: begin  real1=16'b0011110001011011; imag1=16'b0001010101001001;  end  // angle = 0.107910 pi
    12'b000011011110: begin  real1=16'b0011110001010011; imag1=16'b0001010101100000;  end  // angle = 0.108398 pi
    12'b000011011111: begin  real1=16'b0011110001001011; imag1=16'b0001010101111000;  end  // angle = 0.108887 pi
    12'b000011100000: begin  real1=16'b0011110001000010; imag1=16'b0001010110010000;  end  // angle = 0.109375 pi
    12'b000011100001: begin  real1=16'b0011110000111010; imag1=16'b0001010110100111;  end  // angle = 0.109863 pi
    12'b000011100010: begin  real1=16'b0011110000110001; imag1=16'b0001010110111111;  end  // angle = 0.110352 pi
    12'b000011100011: begin  real1=16'b0011110000101001; imag1=16'b0001010111010111;  end  // angle = 0.110840 pi
    12'b000011100100: begin  real1=16'b0011110000100000; imag1=16'b0001010111101110;  end  // angle = 0.111328 pi
    12'b000011100101: begin  real1=16'b0011110000010111; imag1=16'b0001011000000110;  end  // angle = 0.111816 pi
    12'b000011100110: begin  real1=16'b0011110000001111; imag1=16'b0001011000011101;  end  // angle = 0.112305 pi
    12'b000011100111: begin  real1=16'b0011110000000110; imag1=16'b0001011000110101;  end  // angle = 0.112793 pi
    12'b000011101000: begin  real1=16'b0011101111111101; imag1=16'b0001011001001100;  end  // angle = 0.113281 pi
    12'b000011101001: begin  real1=16'b0011101111110101; imag1=16'b0001011001100100;  end  // angle = 0.113770 pi
    12'b000011101010: begin  real1=16'b0011101111101100; imag1=16'b0001011001111100;  end  // angle = 0.114258 pi
    12'b000011101011: begin  real1=16'b0011101111100011; imag1=16'b0001011010010011;  end  // angle = 0.114746 pi
    12'b000011101100: begin  real1=16'b0011101111011010; imag1=16'b0001011010101011;  end  // angle = 0.115234 pi
    12'b000011101101: begin  real1=16'b0011101111010001; imag1=16'b0001011011000010;  end  // angle = 0.115723 pi
    12'b000011101110: begin  real1=16'b0011101111001000; imag1=16'b0001011011011010;  end  // angle = 0.116211 pi
    12'b000011101111: begin  real1=16'b0011101110111111; imag1=16'b0001011011110001;  end  // angle = 0.116699 pi
    12'b000011110000: begin  real1=16'b0011101110110110; imag1=16'b0001011100001001;  end  // angle = 0.117187 pi
    12'b000011110001: begin  real1=16'b0011101110101101; imag1=16'b0001011100100000;  end  // angle = 0.117676 pi
    12'b000011110010: begin  real1=16'b0011101110100100; imag1=16'b0001011100110111;  end  // angle = 0.118164 pi
    12'b000011110011: begin  real1=16'b0011101110011011; imag1=16'b0001011101001111;  end  // angle = 0.118652 pi
    12'b000011110100: begin  real1=16'b0011101110010010; imag1=16'b0001011101100110;  end  // angle = 0.119141 pi
    12'b000011110101: begin  real1=16'b0011101110001000; imag1=16'b0001011101111110;  end  // angle = 0.119629 pi
    12'b000011110110: begin  real1=16'b0011101101111111; imag1=16'b0001011110010101;  end  // angle = 0.120117 pi
    12'b000011110111: begin  real1=16'b0011101101110110; imag1=16'b0001011110101100;  end  // angle = 0.120605 pi
    12'b000011111000: begin  real1=16'b0011101101101101; imag1=16'b0001011111000100;  end  // angle = 0.121094 pi
    12'b000011111001: begin  real1=16'b0011101101100011; imag1=16'b0001011111011011;  end  // angle = 0.121582 pi
    12'b000011111010: begin  real1=16'b0011101101011010; imag1=16'b0001011111110010;  end  // angle = 0.122070 pi
    12'b000011111011: begin  real1=16'b0011101101010000; imag1=16'b0001100000001010;  end  // angle = 0.122559 pi
    12'b000011111100: begin  real1=16'b0011101101000111; imag1=16'b0001100000100001;  end  // angle = 0.123047 pi
    12'b000011111101: begin  real1=16'b0011101100111110; imag1=16'b0001100000111000;  end  // angle = 0.123535 pi
    12'b000011111110: begin  real1=16'b0011101100110100; imag1=16'b0001100001001111;  end  // angle = 0.124023 pi
    12'b000011111111: begin  real1=16'b0011101100101010; imag1=16'b0001100001100111;  end  // angle = 0.124512 pi
    12'b000100000000: begin  real1=16'b0011101100100001; imag1=16'b0001100001111110;  end  // angle = 0.125000 pi
    12'b000100000001: begin  real1=16'b0011101100010111; imag1=16'b0001100010010101;  end  // angle = 0.125488 pi
    12'b000100000010: begin  real1=16'b0011101100001110; imag1=16'b0001100010101100;  end  // angle = 0.125977 pi
    12'b000100000011: begin  real1=16'b0011101100000100; imag1=16'b0001100011000011;  end  // angle = 0.126465 pi
    12'b000100000100: begin  real1=16'b0011101011111010; imag1=16'b0001100011011011;  end  // angle = 0.126953 pi
    12'b000100000101: begin  real1=16'b0011101011110000; imag1=16'b0001100011110010;  end  // angle = 0.127441 pi
    12'b000100000110: begin  real1=16'b0011101011100110; imag1=16'b0001100100001001;  end  // angle = 0.127930 pi
    12'b000100000111: begin  real1=16'b0011101011011101; imag1=16'b0001100100100000;  end  // angle = 0.128418 pi
    12'b000100001000: begin  real1=16'b0011101011010011; imag1=16'b0001100100110111;  end  // angle = 0.128906 pi
    12'b000100001001: begin  real1=16'b0011101011001001; imag1=16'b0001100101001110;  end  // angle = 0.129395 pi
    12'b000100001010: begin  real1=16'b0011101010111111; imag1=16'b0001100101100101;  end  // angle = 0.129883 pi
    12'b000100001011: begin  real1=16'b0011101010110101; imag1=16'b0001100101111100;  end  // angle = 0.130371 pi
    12'b000100001100: begin  real1=16'b0011101010101011; imag1=16'b0001100110010011;  end  // angle = 0.130859 pi
    12'b000100001101: begin  real1=16'b0011101010100001; imag1=16'b0001100110101010;  end  // angle = 0.131348 pi
    12'b000100001110: begin  real1=16'b0011101010010111; imag1=16'b0001100111000001;  end  // angle = 0.131836 pi
    12'b000100001111: begin  real1=16'b0011101010001101; imag1=16'b0001100111011000;  end  // angle = 0.132324 pi
    12'b000100010000: begin  real1=16'b0011101010000010; imag1=16'b0001100111101111;  end  // angle = 0.132812 pi
    12'b000100010001: begin  real1=16'b0011101001111000; imag1=16'b0001101000000110;  end  // angle = 0.133301 pi
    12'b000100010010: begin  real1=16'b0011101001101110; imag1=16'b0001101000011101;  end  // angle = 0.133789 pi
    12'b000100010011: begin  real1=16'b0011101001100100; imag1=16'b0001101000110100;  end  // angle = 0.134277 pi
    12'b000100010100: begin  real1=16'b0011101001011001; imag1=16'b0001101001001011;  end  // angle = 0.134766 pi
    12'b000100010101: begin  real1=16'b0011101001001111; imag1=16'b0001101001100010;  end  // angle = 0.135254 pi
    12'b000100010110: begin  real1=16'b0011101001000101; imag1=16'b0001101001111001;  end  // angle = 0.135742 pi
    12'b000100010111: begin  real1=16'b0011101000111010; imag1=16'b0001101010010000;  end  // angle = 0.136230 pi
    12'b000100011000: begin  real1=16'b0011101000110000; imag1=16'b0001101010100111;  end  // angle = 0.136719 pi
    12'b000100011001: begin  real1=16'b0011101000100101; imag1=16'b0001101010111110;  end  // angle = 0.137207 pi
    12'b000100011010: begin  real1=16'b0011101000011011; imag1=16'b0001101011010100;  end  // angle = 0.137695 pi
    12'b000100011011: begin  real1=16'b0011101000010000; imag1=16'b0001101011101011;  end  // angle = 0.138184 pi
    12'b000100011100: begin  real1=16'b0011101000000110; imag1=16'b0001101100000010;  end  // angle = 0.138672 pi
    12'b000100011101: begin  real1=16'b0011100111111011; imag1=16'b0001101100011001;  end  // angle = 0.139160 pi
    12'b000100011110: begin  real1=16'b0011100111110000; imag1=16'b0001101100110000;  end  // angle = 0.139648 pi
    12'b000100011111: begin  real1=16'b0011100111100110; imag1=16'b0001101101000110;  end  // angle = 0.140137 pi
    12'b000100100000: begin  real1=16'b0011100111011011; imag1=16'b0001101101011101;  end  // angle = 0.140625 pi
    12'b000100100001: begin  real1=16'b0011100111010000; imag1=16'b0001101101110100;  end  // angle = 0.141113 pi
    12'b000100100010: begin  real1=16'b0011100111000101; imag1=16'b0001101110001010;  end  // angle = 0.141602 pi
    12'b000100100011: begin  real1=16'b0011100110111011; imag1=16'b0001101110100001;  end  // angle = 0.142090 pi
    12'b000100100100: begin  real1=16'b0011100110110000; imag1=16'b0001101110111000;  end  // angle = 0.142578 pi
    12'b000100100101: begin  real1=16'b0011100110100101; imag1=16'b0001101111001110;  end  // angle = 0.143066 pi
    12'b000100100110: begin  real1=16'b0011100110011010; imag1=16'b0001101111100101;  end  // angle = 0.143555 pi
    12'b000100100111: begin  real1=16'b0011100110001111; imag1=16'b0001101111111100;  end  // angle = 0.144043 pi
    12'b000100101000: begin  real1=16'b0011100110000100; imag1=16'b0001110000010010;  end  // angle = 0.144531 pi
    12'b000100101001: begin  real1=16'b0011100101111001; imag1=16'b0001110000101001;  end  // angle = 0.145020 pi
    12'b000100101010: begin  real1=16'b0011100101101110; imag1=16'b0001110000111111;  end  // angle = 0.145508 pi
    12'b000100101011: begin  real1=16'b0011100101100011; imag1=16'b0001110001010110;  end  // angle = 0.145996 pi
    12'b000100101100: begin  real1=16'b0011100101011000; imag1=16'b0001110001101100;  end  // angle = 0.146484 pi
    12'b000100101101: begin  real1=16'b0011100101001100; imag1=16'b0001110010000011;  end  // angle = 0.146973 pi
    12'b000100101110: begin  real1=16'b0011100101000001; imag1=16'b0001110010011001;  end  // angle = 0.147461 pi
    12'b000100101111: begin  real1=16'b0011100100110110; imag1=16'b0001110010110000;  end  // angle = 0.147949 pi
    12'b000100110000: begin  real1=16'b0011100100101011; imag1=16'b0001110011000110;  end  // angle = 0.148438 pi
    12'b000100110001: begin  real1=16'b0011100100011111; imag1=16'b0001110011011101;  end  // angle = 0.148926 pi
    12'b000100110010: begin  real1=16'b0011100100010100; imag1=16'b0001110011110011;  end  // angle = 0.149414 pi
    12'b000100110011: begin  real1=16'b0011100100001001; imag1=16'b0001110100001010;  end  // angle = 0.149902 pi
    12'b000100110100: begin  real1=16'b0011100011111101; imag1=16'b0001110100100000;  end  // angle = 0.150391 pi
    12'b000100110101: begin  real1=16'b0011100011110010; imag1=16'b0001110100110110;  end  // angle = 0.150879 pi
    12'b000100110110: begin  real1=16'b0011100011100110; imag1=16'b0001110101001101;  end  // angle = 0.151367 pi
    12'b000100110111: begin  real1=16'b0011100011011011; imag1=16'b0001110101100011;  end  // angle = 0.151855 pi
    12'b000100111000: begin  real1=16'b0011100011001111; imag1=16'b0001110101111001;  end  // angle = 0.152344 pi
    12'b000100111001: begin  real1=16'b0011100011000011; imag1=16'b0001110110010000;  end  // angle = 0.152832 pi
    12'b000100111010: begin  real1=16'b0011100010111000; imag1=16'b0001110110100110;  end  // angle = 0.153320 pi
    12'b000100111011: begin  real1=16'b0011100010101100; imag1=16'b0001110110111100;  end  // angle = 0.153809 pi
    12'b000100111100: begin  real1=16'b0011100010100001; imag1=16'b0001110111010011;  end  // angle = 0.154297 pi
    12'b000100111101: begin  real1=16'b0011100010010101; imag1=16'b0001110111101001;  end  // angle = 0.154785 pi
    12'b000100111110: begin  real1=16'b0011100010001001; imag1=16'b0001110111111111;  end  // angle = 0.155273 pi
    12'b000100111111: begin  real1=16'b0011100001111101; imag1=16'b0001111000010101;  end  // angle = 0.155762 pi
    12'b000101000000: begin  real1=16'b0011100001110001; imag1=16'b0001111000101011;  end  // angle = 0.156250 pi
    12'b000101000001: begin  real1=16'b0011100001100110; imag1=16'b0001111001000010;  end  // angle = 0.156738 pi
    12'b000101000010: begin  real1=16'b0011100001011010; imag1=16'b0001111001011000;  end  // angle = 0.157227 pi
    12'b000101000011: begin  real1=16'b0011100001001110; imag1=16'b0001111001101110;  end  // angle = 0.157715 pi
    12'b000101000100: begin  real1=16'b0011100001000010; imag1=16'b0001111010000100;  end  // angle = 0.158203 pi
    12'b000101000101: begin  real1=16'b0011100000110110; imag1=16'b0001111010011010;  end  // angle = 0.158691 pi
    12'b000101000110: begin  real1=16'b0011100000101010; imag1=16'b0001111010110000;  end  // angle = 0.159180 pi
    12'b000101000111: begin  real1=16'b0011100000011110; imag1=16'b0001111011000110;  end  // angle = 0.159668 pi
    12'b000101001000: begin  real1=16'b0011100000010010; imag1=16'b0001111011011100;  end  // angle = 0.160156 pi
    12'b000101001001: begin  real1=16'b0011100000000101; imag1=16'b0001111011110010;  end  // angle = 0.160645 pi
    12'b000101001010: begin  real1=16'b0011011111111001; imag1=16'b0001111100001000;  end  // angle = 0.161133 pi
    12'b000101001011: begin  real1=16'b0011011111101101; imag1=16'b0001111100011110;  end  // angle = 0.161621 pi
    12'b000101001100: begin  real1=16'b0011011111100001; imag1=16'b0001111100110100;  end  // angle = 0.162109 pi
    12'b000101001101: begin  real1=16'b0011011111010101; imag1=16'b0001111101001010;  end  // angle = 0.162598 pi
    12'b000101001110: begin  real1=16'b0011011111001000; imag1=16'b0001111101100000;  end  // angle = 0.163086 pi
    12'b000101001111: begin  real1=16'b0011011110111100; imag1=16'b0001111101110110;  end  // angle = 0.163574 pi
    12'b000101010000: begin  real1=16'b0011011110110000; imag1=16'b0001111110001100;  end  // angle = 0.164062 pi
    12'b000101010001: begin  real1=16'b0011011110100011; imag1=16'b0001111110100010;  end  // angle = 0.164551 pi
    12'b000101010010: begin  real1=16'b0011011110010111; imag1=16'b0001111110110111;  end  // angle = 0.165039 pi
    12'b000101010011: begin  real1=16'b0011011110001010; imag1=16'b0001111111001101;  end  // angle = 0.165527 pi
    12'b000101010100: begin  real1=16'b0011011101111110; imag1=16'b0001111111100011;  end  // angle = 0.166016 pi
    12'b000101010101: begin  real1=16'b0011011101110001; imag1=16'b0001111111111001;  end  // angle = 0.166504 pi
    12'b000101010110: begin  real1=16'b0011011101100101; imag1=16'b0010000000001111;  end  // angle = 0.166992 pi
    12'b000101010111: begin  real1=16'b0011011101011000; imag1=16'b0010000000100100;  end  // angle = 0.167480 pi
    12'b000101011000: begin  real1=16'b0011011101001011; imag1=16'b0010000000111010;  end  // angle = 0.167969 pi
    12'b000101011001: begin  real1=16'b0011011100111111; imag1=16'b0010000001010000;  end  // angle = 0.168457 pi
    12'b000101011010: begin  real1=16'b0011011100110010; imag1=16'b0010000001100101;  end  // angle = 0.168945 pi
    12'b000101011011: begin  real1=16'b0011011100100101; imag1=16'b0010000001111011;  end  // angle = 0.169434 pi
    12'b000101011100: begin  real1=16'b0011011100011000; imag1=16'b0010000010010001;  end  // angle = 0.169922 pi
    12'b000101011101: begin  real1=16'b0011011100001100; imag1=16'b0010000010100110;  end  // angle = 0.170410 pi
    12'b000101011110: begin  real1=16'b0011011011111111; imag1=16'b0010000010111100;  end  // angle = 0.170898 pi
    12'b000101011111: begin  real1=16'b0011011011110010; imag1=16'b0010000011010001;  end  // angle = 0.171387 pi
    12'b000101100000: begin  real1=16'b0011011011100101; imag1=16'b0010000011100111;  end  // angle = 0.171875 pi
    12'b000101100001: begin  real1=16'b0011011011011000; imag1=16'b0010000011111101;  end  // angle = 0.172363 pi
    12'b000101100010: begin  real1=16'b0011011011001011; imag1=16'b0010000100010010;  end  // angle = 0.172852 pi
    12'b000101100011: begin  real1=16'b0011011010111110; imag1=16'b0010000100101000;  end  // angle = 0.173340 pi
    12'b000101100100: begin  real1=16'b0011011010110001; imag1=16'b0010000100111101;  end  // angle = 0.173828 pi
    12'b000101100101: begin  real1=16'b0011011010100100; imag1=16'b0010000101010011;  end  // angle = 0.174316 pi
    12'b000101100110: begin  real1=16'b0011011010010111; imag1=16'b0010000101101000;  end  // angle = 0.174805 pi
    12'b000101100111: begin  real1=16'b0011011010001010; imag1=16'b0010000101111101;  end  // angle = 0.175293 pi
    12'b000101101000: begin  real1=16'b0011011001111101; imag1=16'b0010000110010011;  end  // angle = 0.175781 pi
    12'b000101101001: begin  real1=16'b0011011001101111; imag1=16'b0010000110101000;  end  // angle = 0.176270 pi
    12'b000101101010: begin  real1=16'b0011011001100010; imag1=16'b0010000110111110;  end  // angle = 0.176758 pi
    12'b000101101011: begin  real1=16'b0011011001010101; imag1=16'b0010000111010011;  end  // angle = 0.177246 pi
    12'b000101101100: begin  real1=16'b0011011001001000; imag1=16'b0010000111101000;  end  // angle = 0.177734 pi
    12'b000101101101: begin  real1=16'b0011011000111010; imag1=16'b0010000111111110;  end  // angle = 0.178223 pi
    12'b000101101110: begin  real1=16'b0011011000101101; imag1=16'b0010001000010011;  end  // angle = 0.178711 pi
    12'b000101101111: begin  real1=16'b0011011000100000; imag1=16'b0010001000101000;  end  // angle = 0.179199 pi
    12'b000101110000: begin  real1=16'b0011011000010010; imag1=16'b0010001000111101;  end  // angle = 0.179688 pi
    12'b000101110001: begin  real1=16'b0011011000000101; imag1=16'b0010001001010011;  end  // angle = 0.180176 pi
    12'b000101110010: begin  real1=16'b0011010111110111; imag1=16'b0010001001101000;  end  // angle = 0.180664 pi
    12'b000101110011: begin  real1=16'b0011010111101010; imag1=16'b0010001001111101;  end  // angle = 0.181152 pi
    12'b000101110100: begin  real1=16'b0011010111011100; imag1=16'b0010001010010010;  end  // angle = 0.181641 pi
    12'b000101110101: begin  real1=16'b0011010111001110; imag1=16'b0010001010100111;  end  // angle = 0.182129 pi
    12'b000101110110: begin  real1=16'b0011010111000001; imag1=16'b0010001010111100;  end  // angle = 0.182617 pi
    12'b000101110111: begin  real1=16'b0011010110110011; imag1=16'b0010001011010010;  end  // angle = 0.183105 pi
    12'b000101111000: begin  real1=16'b0011010110100101; imag1=16'b0010001011100111;  end  // angle = 0.183594 pi
    12'b000101111001: begin  real1=16'b0011010110011000; imag1=16'b0010001011111100;  end  // angle = 0.184082 pi
    12'b000101111010: begin  real1=16'b0011010110001010; imag1=16'b0010001100010001;  end  // angle = 0.184570 pi
    12'b000101111011: begin  real1=16'b0011010101111100; imag1=16'b0010001100100110;  end  // angle = 0.185059 pi
    12'b000101111100: begin  real1=16'b0011010101101110; imag1=16'b0010001100111011;  end  // angle = 0.185547 pi
    12'b000101111101: begin  real1=16'b0011010101100001; imag1=16'b0010001101010000;  end  // angle = 0.186035 pi
    12'b000101111110: begin  real1=16'b0011010101010011; imag1=16'b0010001101100101;  end  // angle = 0.186523 pi
    12'b000101111111: begin  real1=16'b0011010101000101; imag1=16'b0010001101111010;  end  // angle = 0.187012 pi
    12'b000110000000: begin  real1=16'b0011010100110111; imag1=16'b0010001110001110;  end  // angle = 0.187500 pi
    12'b000110000001: begin  real1=16'b0011010100101001; imag1=16'b0010001110100011;  end  // angle = 0.187988 pi
    12'b000110000010: begin  real1=16'b0011010100011011; imag1=16'b0010001110111000;  end  // angle = 0.188477 pi
    12'b000110000011: begin  real1=16'b0011010100001101; imag1=16'b0010001111001101;  end  // angle = 0.188965 pi
    12'b000110000100: begin  real1=16'b0011010011111111; imag1=16'b0010001111100010;  end  // angle = 0.189453 pi
    12'b000110000101: begin  real1=16'b0011010011110001; imag1=16'b0010001111110111;  end  // angle = 0.189941 pi
    12'b000110000110: begin  real1=16'b0011010011100010; imag1=16'b0010010000001011;  end  // angle = 0.190430 pi
    12'b000110000111: begin  real1=16'b0011010011010100; imag1=16'b0010010000100000;  end  // angle = 0.190918 pi
    12'b000110001000: begin  real1=16'b0011010011000110; imag1=16'b0010010000110101;  end  // angle = 0.191406 pi
    12'b000110001001: begin  real1=16'b0011010010111000; imag1=16'b0010010001001010;  end  // angle = 0.191895 pi
    12'b000110001010: begin  real1=16'b0011010010101010; imag1=16'b0010010001011110;  end  // angle = 0.192383 pi
    12'b000110001011: begin  real1=16'b0011010010011011; imag1=16'b0010010001110011;  end  // angle = 0.192871 pi
    12'b000110001100: begin  real1=16'b0011010010001101; imag1=16'b0010010010001000;  end  // angle = 0.193359 pi
    12'b000110001101: begin  real1=16'b0011010001111111; imag1=16'b0010010010011100;  end  // angle = 0.193848 pi
    12'b000110001110: begin  real1=16'b0011010001110000; imag1=16'b0010010010110001;  end  // angle = 0.194336 pi
    12'b000110001111: begin  real1=16'b0011010001100010; imag1=16'b0010010011000101;  end  // angle = 0.194824 pi
    12'b000110010000: begin  real1=16'b0011010001010011; imag1=16'b0010010011011010;  end  // angle = 0.195312 pi
    12'b000110010001: begin  real1=16'b0011010001000101; imag1=16'b0010010011101111;  end  // angle = 0.195801 pi
    12'b000110010010: begin  real1=16'b0011010000110110; imag1=16'b0010010100000011;  end  // angle = 0.196289 pi
    12'b000110010011: begin  real1=16'b0011010000101000; imag1=16'b0010010100011000;  end  // angle = 0.196777 pi
    12'b000110010100: begin  real1=16'b0011010000011001; imag1=16'b0010010100101100;  end  // angle = 0.197266 pi
    12'b000110010101: begin  real1=16'b0011010000001011; imag1=16'b0010010101000001;  end  // angle = 0.197754 pi
    12'b000110010110: begin  real1=16'b0011001111111100; imag1=16'b0010010101010101;  end  // angle = 0.198242 pi
    12'b000110010111: begin  real1=16'b0011001111101101; imag1=16'b0010010101101001;  end  // angle = 0.198730 pi
    12'b000110011000: begin  real1=16'b0011001111011111; imag1=16'b0010010101111110;  end  // angle = 0.199219 pi
    12'b000110011001: begin  real1=16'b0011001111010000; imag1=16'b0010010110010010;  end  // angle = 0.199707 pi
    12'b000110011010: begin  real1=16'b0011001111000001; imag1=16'b0010010110100110;  end  // angle = 0.200195 pi
    12'b000110011011: begin  real1=16'b0011001110110010; imag1=16'b0010010110111011;  end  // angle = 0.200684 pi
    12'b000110011100: begin  real1=16'b0011001110100011; imag1=16'b0010010111001111;  end  // angle = 0.201172 pi
    12'b000110011101: begin  real1=16'b0011001110010101; imag1=16'b0010010111100011;  end  // angle = 0.201660 pi
    12'b000110011110: begin  real1=16'b0011001110000110; imag1=16'b0010010111111000;  end  // angle = 0.202148 pi
    12'b000110011111: begin  real1=16'b0011001101110111; imag1=16'b0010011000001100;  end  // angle = 0.202637 pi
    12'b000110100000: begin  real1=16'b0011001101101000; imag1=16'b0010011000100000;  end  // angle = 0.203125 pi
    12'b000110100001: begin  real1=16'b0011001101011001; imag1=16'b0010011000110100;  end  // angle = 0.203613 pi
    12'b000110100010: begin  real1=16'b0011001101001010; imag1=16'b0010011001001000;  end  // angle = 0.204102 pi
    12'b000110100011: begin  real1=16'b0011001100111011; imag1=16'b0010011001011100;  end  // angle = 0.204590 pi
    12'b000110100100: begin  real1=16'b0011001100101100; imag1=16'b0010011001110001;  end  // angle = 0.205078 pi
    12'b000110100101: begin  real1=16'b0011001100011101; imag1=16'b0010011010000101;  end  // angle = 0.205566 pi
    12'b000110100110: begin  real1=16'b0011001100001101; imag1=16'b0010011010011001;  end  // angle = 0.206055 pi
    12'b000110100111: begin  real1=16'b0011001011111110; imag1=16'b0010011010101101;  end  // angle = 0.206543 pi
    12'b000110101000: begin  real1=16'b0011001011101111; imag1=16'b0010011011000001;  end  // angle = 0.207031 pi
    12'b000110101001: begin  real1=16'b0011001011100000; imag1=16'b0010011011010101;  end  // angle = 0.207520 pi
    12'b000110101010: begin  real1=16'b0011001011010000; imag1=16'b0010011011101001;  end  // angle = 0.208008 pi
    12'b000110101011: begin  real1=16'b0011001011000001; imag1=16'b0010011011111101;  end  // angle = 0.208496 pi
    12'b000110101100: begin  real1=16'b0011001010110010; imag1=16'b0010011100010001;  end  // angle = 0.208984 pi
    12'b000110101101: begin  real1=16'b0011001010100011; imag1=16'b0010011100100100;  end  // angle = 0.209473 pi
    12'b000110101110: begin  real1=16'b0011001010010011; imag1=16'b0010011100111000;  end  // angle = 0.209961 pi
    12'b000110101111: begin  real1=16'b0011001010000100; imag1=16'b0010011101001100;  end  // angle = 0.210449 pi
    12'b000110110000: begin  real1=16'b0011001001110100; imag1=16'b0010011101100000;  end  // angle = 0.210938 pi
    12'b000110110001: begin  real1=16'b0011001001100101; imag1=16'b0010011101110100;  end  // angle = 0.211426 pi
    12'b000110110010: begin  real1=16'b0011001001010101; imag1=16'b0010011110001000;  end  // angle = 0.211914 pi
    12'b000110110011: begin  real1=16'b0011001001000110; imag1=16'b0010011110011011;  end  // angle = 0.212402 pi
    12'b000110110100: begin  real1=16'b0011001000110110; imag1=16'b0010011110101111;  end  // angle = 0.212891 pi
    12'b000110110101: begin  real1=16'b0011001000100111; imag1=16'b0010011111000011;  end  // angle = 0.213379 pi
    12'b000110110110: begin  real1=16'b0011001000010111; imag1=16'b0010011111010110;  end  // angle = 0.213867 pi
    12'b000110110111: begin  real1=16'b0011001000000111; imag1=16'b0010011111101010;  end  // angle = 0.214355 pi
    12'b000110111000: begin  real1=16'b0011000111111000; imag1=16'b0010011111111110;  end  // angle = 0.214844 pi
    12'b000110111001: begin  real1=16'b0011000111101000; imag1=16'b0010100000010001;  end  // angle = 0.215332 pi
    12'b000110111010: begin  real1=16'b0011000111011000; imag1=16'b0010100000100101;  end  // angle = 0.215820 pi
    12'b000110111011: begin  real1=16'b0011000111001000; imag1=16'b0010100000111000;  end  // angle = 0.216309 pi
    12'b000110111100: begin  real1=16'b0011000110111001; imag1=16'b0010100001001100;  end  // angle = 0.216797 pi
    12'b000110111101: begin  real1=16'b0011000110101001; imag1=16'b0010100001100000;  end  // angle = 0.217285 pi
    12'b000110111110: begin  real1=16'b0011000110011001; imag1=16'b0010100001110011;  end  // angle = 0.217773 pi
    12'b000110111111: begin  real1=16'b0011000110001001; imag1=16'b0010100010000110;  end  // angle = 0.218262 pi
    12'b000111000000: begin  real1=16'b0011000101111001; imag1=16'b0010100010011010;  end  // angle = 0.218750 pi
    12'b000111000001: begin  real1=16'b0011000101101001; imag1=16'b0010100010101101;  end  // angle = 0.219238 pi
    12'b000111000010: begin  real1=16'b0011000101011001; imag1=16'b0010100011000001;  end  // angle = 0.219727 pi
    12'b000111000011: begin  real1=16'b0011000101001001; imag1=16'b0010100011010100;  end  // angle = 0.220215 pi
    12'b000111000100: begin  real1=16'b0011000100111001; imag1=16'b0010100011100111;  end  // angle = 0.220703 pi
    12'b000111000101: begin  real1=16'b0011000100101001; imag1=16'b0010100011111011;  end  // angle = 0.221191 pi
    12'b000111000110: begin  real1=16'b0011000100011001; imag1=16'b0010100100001110;  end  // angle = 0.221680 pi
    12'b000111000111: begin  real1=16'b0011000100001001; imag1=16'b0010100100100001;  end  // angle = 0.222168 pi
    12'b000111001000: begin  real1=16'b0011000011111001; imag1=16'b0010100100110101;  end  // angle = 0.222656 pi
    12'b000111001001: begin  real1=16'b0011000011101000; imag1=16'b0010100101001000;  end  // angle = 0.223145 pi
    12'b000111001010: begin  real1=16'b0011000011011000; imag1=16'b0010100101011011;  end  // angle = 0.223633 pi
    12'b000111001011: begin  real1=16'b0011000011001000; imag1=16'b0010100101101110;  end  // angle = 0.224121 pi
    12'b000111001100: begin  real1=16'b0011000010111000; imag1=16'b0010100110000001;  end  // angle = 0.224609 pi
    12'b000111001101: begin  real1=16'b0011000010100111; imag1=16'b0010100110010100;  end  // angle = 0.225098 pi
    12'b000111001110: begin  real1=16'b0011000010010111; imag1=16'b0010100110100111;  end  // angle = 0.225586 pi
    12'b000111001111: begin  real1=16'b0011000010000111; imag1=16'b0010100110111011;  end  // angle = 0.226074 pi
    12'b000111010000: begin  real1=16'b0011000001110110; imag1=16'b0010100111001110;  end  // angle = 0.226562 pi
    12'b000111010001: begin  real1=16'b0011000001100110; imag1=16'b0010100111100001;  end  // angle = 0.227051 pi
    12'b000111010010: begin  real1=16'b0011000001010101; imag1=16'b0010100111110100;  end  // angle = 0.227539 pi
    12'b000111010011: begin  real1=16'b0011000001000101; imag1=16'b0010101000000111;  end  // angle = 0.228027 pi
    12'b000111010100: begin  real1=16'b0011000000110100; imag1=16'b0010101000011010;  end  // angle = 0.228516 pi
    12'b000111010101: begin  real1=16'b0011000000100100; imag1=16'b0010101000101100;  end  // angle = 0.229004 pi
    12'b000111010110: begin  real1=16'b0011000000010011; imag1=16'b0010101000111111;  end  // angle = 0.229492 pi
    12'b000111010111: begin  real1=16'b0011000000000010; imag1=16'b0010101001010010;  end  // angle = 0.229980 pi
    12'b000111011000: begin  real1=16'b0010111111110010; imag1=16'b0010101001100101;  end  // angle = 0.230469 pi
    12'b000111011001: begin  real1=16'b0010111111100001; imag1=16'b0010101001111000;  end  // angle = 0.230957 pi
    12'b000111011010: begin  real1=16'b0010111111010000; imag1=16'b0010101010001011;  end  // angle = 0.231445 pi
    12'b000111011011: begin  real1=16'b0010111111000000; imag1=16'b0010101010011101;  end  // angle = 0.231934 pi
    12'b000111011100: begin  real1=16'b0010111110101111; imag1=16'b0010101010110000;  end  // angle = 0.232422 pi
    12'b000111011101: begin  real1=16'b0010111110011110; imag1=16'b0010101011000011;  end  // angle = 0.232910 pi
    12'b000111011110: begin  real1=16'b0010111110001101; imag1=16'b0010101011010110;  end  // angle = 0.233398 pi
    12'b000111011111: begin  real1=16'b0010111101111101; imag1=16'b0010101011101000;  end  // angle = 0.233887 pi
    12'b000111100000: begin  real1=16'b0010111101101100; imag1=16'b0010101011111011;  end  // angle = 0.234375 pi
    12'b000111100001: begin  real1=16'b0010111101011011; imag1=16'b0010101100001101;  end  // angle = 0.234863 pi
    12'b000111100010: begin  real1=16'b0010111101001010; imag1=16'b0010101100100000;  end  // angle = 0.235352 pi
    12'b000111100011: begin  real1=16'b0010111100111001; imag1=16'b0010101100110011;  end  // angle = 0.235840 pi
    12'b000111100100: begin  real1=16'b0010111100101000; imag1=16'b0010101101000101;  end  // angle = 0.236328 pi
    12'b000111100101: begin  real1=16'b0010111100010111; imag1=16'b0010101101011000;  end  // angle = 0.236816 pi
    12'b000111100110: begin  real1=16'b0010111100000110; imag1=16'b0010101101101010;  end  // angle = 0.237305 pi
    12'b000111100111: begin  real1=16'b0010111011110101; imag1=16'b0010101101111101;  end  // angle = 0.237793 pi
    12'b000111101000: begin  real1=16'b0010111011100100; imag1=16'b0010101110001111;  end  // angle = 0.238281 pi
    12'b000111101001: begin  real1=16'b0010111011010011; imag1=16'b0010101110100001;  end  // angle = 0.238770 pi
    12'b000111101010: begin  real1=16'b0010111011000010; imag1=16'b0010101110110100;  end  // angle = 0.239258 pi
    12'b000111101011: begin  real1=16'b0010111010110000; imag1=16'b0010101111000110;  end  // angle = 0.239746 pi
    12'b000111101100: begin  real1=16'b0010111010011111; imag1=16'b0010101111011000;  end  // angle = 0.240234 pi
    12'b000111101101: begin  real1=16'b0010111010001110; imag1=16'b0010101111101011;  end  // angle = 0.240723 pi
    12'b000111101110: begin  real1=16'b0010111001111101; imag1=16'b0010101111111101;  end  // angle = 0.241211 pi
    12'b000111101111: begin  real1=16'b0010111001101011; imag1=16'b0010110000001111;  end  // angle = 0.241699 pi
    12'b000111110000: begin  real1=16'b0010111001011010; imag1=16'b0010110000100001;  end  // angle = 0.242188 pi
    12'b000111110001: begin  real1=16'b0010111001001001; imag1=16'b0010110000110100;  end  // angle = 0.242676 pi
    12'b000111110010: begin  real1=16'b0010111000110111; imag1=16'b0010110001000110;  end  // angle = 0.243164 pi
    12'b000111110011: begin  real1=16'b0010111000100110; imag1=16'b0010110001011000;  end  // angle = 0.243652 pi
    12'b000111110100: begin  real1=16'b0010111000010101; imag1=16'b0010110001101010;  end  // angle = 0.244141 pi
    12'b000111110101: begin  real1=16'b0010111000000011; imag1=16'b0010110001111100;  end  // angle = 0.244629 pi
    12'b000111110110: begin  real1=16'b0010110111110010; imag1=16'b0010110010001110;  end  // angle = 0.245117 pi
    12'b000111110111: begin  real1=16'b0010110111100000; imag1=16'b0010110010100000;  end  // angle = 0.245605 pi
    12'b000111111000: begin  real1=16'b0010110111001111; imag1=16'b0010110010110010;  end  // angle = 0.246094 pi
    12'b000111111001: begin  real1=16'b0010110110111101; imag1=16'b0010110011000100;  end  // angle = 0.246582 pi
    12'b000111111010: begin  real1=16'b0010110110101011; imag1=16'b0010110011010110;  end  // angle = 0.247070 pi
    12'b000111111011: begin  real1=16'b0010110110011010; imag1=16'b0010110011101000;  end  // angle = 0.247559 pi
    12'b000111111100: begin  real1=16'b0010110110001000; imag1=16'b0010110011111010;  end  // angle = 0.248047 pi
    12'b000111111101: begin  real1=16'b0010110101110110; imag1=16'b0010110100001100;  end  // angle = 0.248535 pi
    12'b000111111110: begin  real1=16'b0010110101100101; imag1=16'b0010110100011110;  end  // angle = 0.249023 pi
    12'b000111111111: begin  real1=16'b0010110101010011; imag1=16'b0010110100101111;  end  // angle = 0.249512 pi
    12'b001000000000: begin  real1=16'b0010110101000001; imag1=16'b0010110101000001;  end  // angle = 0.250000 pi
  endcase
end

endmodule
