
module Top_tb;
reg [3:0] inp1;
reg [3:0] inp2;
reg [3:0] inp3;
reg [3:0] inp4;
reg [3:0] inp5;
reg [3:0] inp6;
wire [5:0] answerp;
Top Toptestbench (inp1 [3:0],inp2 [3:0],inp3 [3:0],inp4 [3:0],inp5 [3:0],inp6 [3:0],answerp [5:0]);

initial 
begin
$monitor ($time, "inp1 = %b \t inp2 = %b \t inp3 = %b \t inp4 = %b \t inp5 = %b \t inp6 = %b \t answerp = %b \t",inp1[3:0],inp2[3:0],inp3[3:0],inp4[3:0],inp5[3:0],inp6[3:0],answerp[5:0]);
#5;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0001;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0001;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0001;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0001;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0001;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0001;
#50;
inp1[3:0] = 4'b1111;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b1111;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b1111;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b1111;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b1111;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b1111;
#50;
inp1[3:0] = 4'b0111; //7
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0111;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0111;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0111;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0111;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0111;
#50;
inp1[3:0] = 4'b1000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b1000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b1000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b1000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b1000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b1000;
#50;
inp1[3:0] = 4'b0001;
inp2[3:0] = 4'b0001;
inp3[3:0] = 4'b0001;
inp4[3:0] = 4'b0001;
inp5[3:0] = 4'b0001;
inp6[3:0] = 4'b0001;
#50;
inp1[3:0] = 4'b1111;
inp2[3:0] = 4'b1111;
inp3[3:0] = 4'b1111;
inp4[3:0] = 4'b1111;
inp5[3:0] = 4'b1111;
inp6[3:0] = 4'b1111;
#50;
inp1[3:0] = 4'b0001;
inp2[3:0] = 4'b0010;
inp3[3:0] = 4'b0011;
inp4[3:0] = 4'b0100;
inp5[3:0] = 4'b0101;
inp6[3:0] = 4'b0110;
#50;
inp1[3:0] = 4'b0110;
inp2[3:0] = 4'b0101;
inp3[3:0] = 4'b0101;
inp4[3:0] = 4'b0101;
inp5[3:0] = 4'b0101;
inp6[3:0] = 4'b0101;
#50;
inp1[3:0] = 4'b0000;
inp2[3:0] = 4'b0000;
inp3[3:0] = 4'b0000;
inp4[3:0] = 4'b0000;
inp5[3:0] = 4'b0000;
inp6[3:0] = 4'b0000;
#50;
inp1[3:0] = 4'b1001; //-7
inp2[3:0] = 4'b1011; //-5
inp3[3:0] = 4'b1011; //-5
inp4[3:0] = 4'b1011; //-5
inp5[3:0] = 4'b1011; //-5
inp6[3:0] = 4'b1011; //-5
#100;
end
endmodule
