module Inverter2 (in,out);
input in;
output out;
assign out = ~in;
endmodule;
