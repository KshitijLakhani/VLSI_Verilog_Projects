// Trial verilog code for implementing inverter
module Inverter (in,out);

input in;
output out;

assign out = ~ in;
endmodule
