module Top (
input [7:0] multiplicand,
input [7:0] multiplier,
output reg [15:0] answer,
output reg [15:0] answer_temp);
wire [15:0] pp0;
wire [15:0] pp1;
wire [15:0] pp2;
wire [15:0] pp3;
wire [15:0] pp4;
wire [15:0] pp5;
wire [15:0] pp6;
wire [15:0] pp7;

wire [15:0] stage1_line1;
wire [15:0] stage1_line2;
wire [15:0] stage2_line1;
wire [15:0] stage2_line2;

wire [15:0] stage3_line1;
wire [15:0] stage3_line2;

wire multiplicand_negative;
wire multiplier_negative;
wire maxneg_multiplier;
wire maxneg_multiplicand;

//reg [15:0] answer_temp;

//wire [15:0] temp;

partial_product_generator mod1(multiplicand[7:0],multiplier[7:0],pp0[15:0],pp1[15:0],pp2[15:0],pp3[15:0],pp4[15:0],pp5[15:0],pp6[15:0],pp7[15:0],multiplicand_negative,multiplier_negative,maxneg_multiplicand,maxneg_multiplier);
stage1 mod2(pp0[15:0],pp1[15:0],pp2[15:0],pp3[15:0],stage1_line1[15:0],stage1_line2[15:0]);
stage2 mod3(pp4[15:0],pp5[15:0],pp6[15:0],pp7[15:0],stage2_line1[15:0],stage2_line2[15:0]);
stage3 mod4(stage1_line1[15:0],stage1_line2[15:0],stage2_line1[15:0],stage2_line2[15:0],stage3_line1[15:0],stage3_line2[15:0]);



always @(*)
begin
answer_temp[15:0]=stage3_line1[15:0] + stage3_line2[15:0] + {5'b00000,4'b1111,7'b0000000};

if((multiplicand_negative ^ multiplier_negative)==1)
begin
answer[15:0]=(~answer_temp[15:0]) + 15'b00000001;
/*if (maxneg_multiplier==1)
begin
answer[15:0]=(~answer_temp[15:0]) + 8'b00000001 + {};
end
if(maxneg_multiplicand==1)
begin
answer[15:0]=(~(answer_temp[15:0] + {8'b00000000,multiplier[7:0]})) + 8'b00000001;
end*/

end

else 
begin
/*if((maxneg_multiplier==1) & (maxneg_multiplicand==1))
begin
answer[15:0]=answer_temp[15:0] + 16'b0000000011111111;
end
else
begin
answer[15:0]=answer_temp[15:0];
end*/
answer[15:0]=answer_temp[15:0];
end
end
endmodule

module stage1 (
input [15:0] pp0,
input [15:0] pp1,
input [15:0] pp2,
input [15:0] pp3,
output [15:0] stage1_line1,
output [15:0] stage1_line2);

assign stage1_line2[15:12]=4'b1110;  //brick wall ensures that MSBs 11 from 1111100 gets thrown off
assign stage1_line1[15:12]=4'b0000;

assign stage1_line1[1:0]={pp0[1],pp0[0]};
assign stage1_line2[2:0]={1'b0,pp1[1],1'b0};

wire cs0_c0,cs1_c0,cs2_c0,cs3_c0,cs4_c0,cs5_c0,cs6_c0,cs7_c0;
//instantiation of 9 4is2 carry save adder
carrysave_4is2 cs0({pp0[2],pp1[2],pp2[2],2'b00},cs0_c0,stage1_line2[3],stage1_line1[2]);
carrysave_4is2 cs1({pp0[3],pp1[3],pp2[3],pp3[3],cs0_c0},cs1_c0,stage1_line2[4],stage1_line1[3]);
carrysave_4is2 cs2({pp0[4],pp1[4],pp2[4],pp3[4],cs1_c0},cs2_c0,stage1_line2[5],stage1_line1[4]);
carrysave_4is2 cs3({pp0[5],pp1[5],pp2[5],pp3[5],cs2_c0},cs3_c0,stage1_line2[6],stage1_line1[5]);
carrysave_4is2 cs4({pp0[6],pp1[6],pp2[6],pp3[6],cs3_c0},cs4_c0,stage1_line2[7],stage1_line1[6]);
carrysave_4is2 cs5({~pp0[7],pp1[7],pp2[7],pp3[7],cs4_c0},cs5_c0,stage1_line2[8],stage1_line1[7]);
carrysave_4is2 cs6({1'b1,~pp1[8],pp2[8],pp3[8],cs5_c0},cs6_c0,stage1_line2[9],stage1_line1[8]);
carrysave_4is2 cs7({1'b1,1'b1,~pp2[9],pp3[9],cs6_c0},cs7_c0,stage1_line2[10],stage1_line1[9]);
carrysave_4is2 cs8({1'b1,1'b1,1'b1,~pp3[10],cs7_c0},stage1_line1[11],stage1_line2[11],stage1_line1[10]);
//Accomodate for the extra 1's

endmodule

module stage2 (
input [15:0] pp4,
input [15:0] pp5,
input [15:0] pp6,
input [15:0] pp7,
output [15:0] stage2_line1,
output [15:0] stage2_line2);

assign stage2_line1[5:0]={pp4[5],pp4[4],4'b0000};
assign stage2_line2[6:0]={1'b0,pp5[5],5'b00000};

wire cs9_c0,cs10_c0,cs11_c0,cs12_c0,cs13_c0,cs14_c0,cs15_c0,cs16_c0,cs17_c0;

carrysave_4is2 cs9({pp4[6],pp5[6],pp6[6],2'b00},cs9_c0,stage2_line2[7],stage2_line1[6]);
carrysave_4is2 cs10({pp4[7],pp5[7],pp6[7],pp7[7],cs9_c0},cs10_c0,stage2_line2[8],stage2_line1[7]);
carrysave_4is2 cs11({pp4[8],pp5[8],pp6[8],pp7[8],cs10_c0},cs11_c0,stage2_line2[9],stage2_line1[8]);
carrysave_4is2 cs12({pp4[9],pp5[9],pp6[9],pp7[9],cs11_c0},cs12_c0,stage2_line2[10],stage2_line1[9]);
carrysave_4is2 cs13({pp4[10],pp5[10],pp6[10],pp7[10],cs12_c0},cs13_c0,stage2_line2[11],stage2_line1[10]);
carrysave_4is2 cs14({pp4[11],pp5[11],pp6[11],pp7[11],cs13_c0},cs14_c0,stage2_line2[12],stage2_line1[11]);
carrysave_4is2 cs15({pp4[12],pp5[12],pp6[12],pp7[12],cs14_c0},cs15_c0,stage2_line2[13],stage2_line1[12]);
carrysave_4is2 cs16({pp4[13],pp5[13],pp6[13],pp7[13],cs15_c0},cs16_c0,stage2_line2[14],stage2_line1[13]);
carrysave_4is2 cs17({pp4[14],pp5[14],pp6[14],pp7[14],cs16_c0},cs17_c0,stage2_line2[15],stage2_line1[14]);
carrysave_4is2 cs18({pp4[15],pp5[15],pp6[15],pp7[15],cs17_c0}, , ,stage2_line1[15]);

endmodule

module stage3 (
input [15:0] stage1_line1,
input [15:0] stage1_line2,
input [15:0] stage2_line1,
input [15:0] stage2_line2,
output [15:0] stage3_line1,
output [15:0] stage3_line2);

assign stage3_line2[0]=1'b0;

carrysave_4is2 cs19({stage1_line1[0],stage1_line2[0],stage2_line1[0],stage2_line2[0],1'b0},cs19_c0,stage3_line2[1],stage3_line1[0]);
carrysave_4is2 cs20({stage1_line1[1],stage1_line2[1],stage2_line1[1],stage2_line2[1],cs19_c0},cs20_c0,stage3_line2[2],stage3_line1[1]);
carrysave_4is2 cs21({stage1_line1[2],stage1_line2[2],stage2_line1[2],stage2_line2[2],cs20_c0},cs21_c0,stage3_line2[3],stage3_line1[2]);
carrysave_4is2 cs22({stage1_line1[3],stage1_line2[3],stage2_line1[3],stage2_line2[3],cs21_c0},cs22_c0,stage3_line2[4],stage3_line1[3]);
carrysave_4is2 cs23({stage1_line1[4],stage1_line2[4],stage2_line1[4],stage2_line2[4],cs22_c0},cs23_c0,stage3_line2[5],stage3_line1[4]);
carrysave_4is2 cs24({stage1_line1[5],stage1_line2[5],stage2_line1[5],stage2_line2[5],cs23_c0},cs24_c0,stage3_line2[6],stage3_line1[5]);
carrysave_4is2 cs25({stage1_line1[6],stage1_line2[6],stage2_line1[6],stage2_line2[6],cs24_c0},cs25_c0,stage3_line2[7],stage3_line1[6]);
carrysave_4is2 cs26({stage1_line1[7],stage1_line2[7],stage2_line1[7],stage2_line2[7],cs25_c0},cs26_c0,stage3_line2[8],stage3_line1[7]);
carrysave_4is2 cs27({stage1_line1[8],stage1_line2[8],stage2_line1[8],stage2_line2[8],cs26_c0},cs27_c0,stage3_line2[9],stage3_line1[8]);
carrysave_4is2 cs28({stage1_line1[9],stage1_line2[9],stage2_line1[9],stage2_line2[9],cs27_c0},cs28_c0,stage3_line2[10],stage3_line1[9]);
carrysave_4is2 cs29({stage1_line1[10],stage1_line2[10],stage2_line1[10],stage2_line2[10],cs28_c0},cs29_c0,stage3_line2[11],stage3_line1[10]);
carrysave_4is2 cs30({stage1_line1[11],stage1_line2[11],stage2_line1[11],stage2_line2[11],cs29_c0},cs30_c0,stage3_line2[12],stage3_line1[11]);
carrysave_4is2 cs31({stage1_line1[12],stage1_line2[12],stage2_line1[12],stage2_line2[12],cs30_c0},cs31_c0,stage3_line2[13],stage3_line1[12]);
carrysave_4is2 cs32({stage1_line1[13],stage1_line2[13],stage2_line1[13],stage2_line2[13],cs31_c0},cs32_c0,stage3_line2[14],stage3_line1[13]);
carrysave_4is2 cs33({stage1_line1[14],stage1_line2[14],stage2_line1[14],stage2_line2[14],cs32_c0},cs33_c0,stage3_line2[15],stage3_line1[14]);
carrysave_4is2 cs34({stage1_line1[15],stage1_line2[15],stage2_line1[15],stage2_line2[15],cs33_c0}, , ,stage3_line1[15]);
endmodule

module partial_product_generator(
input reg [7:0] multiplicand,
input reg [7:0] multiplier,
output reg [15:0] pp0,
output reg [15:0] pp1,
output reg [15:0] pp2,
output reg [15:0] pp3,
output reg [15:0] pp4,
output reg [15:0] pp5,
output reg [15:0] pp6,
output reg [15:0] pp7,
output reg plicand_negative,
output reg plier_negative,
output reg flag_maxneg_multiplicand,
output reg flag_maxneg_multiplier);

reg [7:0] plier;
reg [7:0] plicand;
//reg [7:0] temp
always @(*)
begin
//code for negative inputs
plier_negative=1'b0;
plicand_negative=1'b0;
flag_maxneg_multiplier=1'b0;
flag_maxneg_multiplicand=1'b0;

plier[7:0]=multiplier[7:0];
plicand[7:0]=multiplicand[7:0];

if (multiplier[7]==1)
begin
plier[7:0]= (~ multiplier[7:0]) + (8'b00000001);
plier_negative=1'b1;
if (multiplier[7:0] == 8'b10000000)
begin
flag_maxneg_multiplier=1'b1;
end
end

if (plier[0]==0)
begin
pp0[15:0]=16'h0000;
end
else
begin
pp0[15:0]={plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7:0]};
if (multiplicand[7:0] == 8'b10000000)
begin
pp0[15:0]={8'b00000000,plicand[7:0]};
end
end


if (multiplicand[7]==1)
begin
plicand[7:0]= (~ multiplicand[7:0]) + (8'b00000001);
plicand_negative=1'b1;
if (multiplicand[7:0] == 8'b10000000)
begin
flag_maxneg_multiplicand=1'b1;
//temp[7:0]=multiplicand[7:0]
end
end

if (plier[1]==0)
begin
pp1[15:0]=16'h0000;
end
else
begin
pp1[15:0]={plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7:0],1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp1[15:0]={7'b0000000,plicand[7:0],1'b0};
end
end

if (plier[2]==0)
begin
pp2[15:0]=16'h0000;
end
else
begin
pp2[15:0]={plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7:0],1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp2[15:0]={6'b000000,plicand[7:0],2'b00};
end
end

if (plier[3]==0)
begin
pp3[15:0]=16'h0000;
end
else
begin
pp3[15:0]={plicand[7],plicand[7],plicand[7],plicand[7],plicand[7],plicand[7:0],1'b0,1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp3[15:0]={5'b00000,plicand[7:0],3'b000};
end
end

if (plier[4]==0)
begin
pp4[15:0]=16'h0000;
end
else
begin
pp4[15:0]={plicand[7],plicand[7],plicand[7],plicand[7],plicand[7:0],1'b0,1'b0,1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp4[15:0]={4'b0000,plicand[7:0],4'b0000};
end
end

if (plier[5]==0)
begin
pp5[15:0]=16'h0000;
end
else
begin
pp5[15:0]={plicand[7],plicand[7],plicand[7],plicand[7:0],1'b0,1'b0,1'b0,1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp5[15:0]={3'b000,plicand[7:0],5'b00000};
end
end

if (plier[6]==0)
begin
pp6[15:0]=16'h0000;
end
else
begin
pp6[15:0]={plicand[7],plicand[7],plicand[7:0],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp6[15:0]={2'b00,plicand[7:0],6'b000000};
end
end

if (plier[7]==0)
begin
pp7[15:0]=16'h0000;
end
else
begin
pp7[15:0]={plicand[7],plicand[7:0],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
if (multiplicand[7:0] == 8'b10000000)
begin
pp7[15:0]={1'b0,plicand[7:0],7'b0000000};
end
end
end

endmodule
module carrysave_4is2 (
input [4:0] in,
output c0,
output c1,
output sum
);
wire connection;
FullAdder FA0 (in[4],in[3],in[2],connection,c0);
FullAdder FA1 (connection,in[1],in[0],sum,c1);
endmodule

module FullAdder(
input in1,
input in2,
input cin,
output sum,
output cout
);
assign sum = (in1 ^ in2) ^ cin;
assign cout = (in1 & in2) | (cin & (in1 ^ in2));
endmodule
