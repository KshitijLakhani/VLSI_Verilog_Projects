module Top_tb;
reg [4:0] a;
reg [4:0] b;
reg [4:0] c;
wire [8:0] addition;

Top testbench_adddition (a[4:0],b[4:0],c[4:0],addition[8:0]);

initial
begin
$monitor ($time,"a = %b \t b = %b \t c = %b \t addition = %b \n",a[4:0],b[4:0],c[4:0],addition[8:0]);
#10
a[4:0] = 10000;
b[4:0] = 10000;
c[4:0] = 01111;
#50;
a[4:0] = 10010;
b[4:0] = 10100;
c[4:0] = 11111;
#50;
a[4:0] = 10101;
b[4:0] = 10001;
c[4:0] = 01011;
#50;
a[4:0] = 10110;
b[4:0] = 11100;
c[4:0] = 11011;
#50;
a[4:0] = 00000;
b[4:0] = 00000;
c[4:0] = 00000;
#50;
a[4:0] = 11111;
b[4:0] = 11111;
c[4:0] = 11111;
#50;
a[4:0] = 10000;
b[4:0] = 1000;
c[4:0] = 10011;
#50;
a[4:0] = 00111;
b[4:0] = 11100;
c[4:0] = 11111;
#50;
a[4:0] = 01100;
b[4:0] = 01100;
c[4:0] = 01111;
#50;
a[4:0] = 00111;
b[4:0] = 00101;
c[4:0] = 01001;
#50;
a[4:0] = 10101;
b[4:0] = 10101;
c[4:0] = 11010;
#50;
a[4:0] = 00001;
b[4:0] = 00001;
c[4:0] = 00001;
#50;
a[4:0] = 00100;
b[4:0] = 00100;
c[4:0] = 01100;
#50;
a[4:0] = 11011;
b[4:0] = 11011;
c[4:0] = 11011;
#50;
a[4:0] = 01110;
b[4:0] = 00001;
c[4:0] = 00101;
#50;
a[4:0] = 00111;
b[4:0] = 10100;
c[4:0] = 01011;
#50;
end
endmodule
